["Voluptatum quam sunt et odio aut voluptas. Sit eum aspernatur quo deleniti a consequuntur autem. Accusantium occaecati consequatur est nihil veritatis. Autem omnis ea ut. Sit ipsum vel inventore minus.", "In placeat culpa ratione autem dolores dolor. Autem nemo maxime ducimus quis corrupti. Iusto nisi neque incidunt eos.", "Nemo ea aut autem nesciunt quia tenetur. Cupiditate quam provident tempore aspernatur et est. Dignissimos aut rerum maiores.", "Placeat nihil nostrum consectetur minima fugiat sit. Consequatur molestiae tempore est eum. Provident ratione nobis amet totam.", "Optio magnam sint eveniet vero fugiat nihil. Eveniet cum vel debitis nihil nemo ipsum fuga. Quaerat quidem veniam sit tempora numquam dolorem. Sapiente nostrum doloremque. Doloribus omnis sed non veritatis minus et dolorem."]