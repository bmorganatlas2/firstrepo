["Officia quae quis temporibus at. Laudantium dolores in. Ullam soluta sit aliquam odit illum repellendus. Et sit ratione eum asperiores quia numquam.", "Non possimus maxime dolorem eos error facilis voluptas. Necessitatibus debitis voluptatem omnis commodi aliquid. Molestias dolore ipsa neque consequuntur et ipsam. Soluta fugit optio est quas eum nisi.", "Ex et a. Nesciunt aut et nobis. Doloremque inventore rerum rem. Saepe eveniet sed dolore impedit inventore enim voluptatibus. Non cupiditate porro.", "Dolorum culpa deserunt accusantium. Delectus impedit necessitatibus officiis numquam quos incidunt repellendus. Rerum et qui eveniet. Aut consequatur commodi autem totam voluptatem animi laboriosam."]