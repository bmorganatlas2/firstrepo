["Est earum quam eligendi explicabo ipsa est. Optio a eaque provident quos rem consequatur. Nam qui officiis vel illo eaque qui. Voluptatem fugiat molestiae natus ea cupiditate iure.", "Adipisci alias quis velit. Autem est ut omnis mollitia numquam fugiat. Laborum sed nisi quidem excepturi et et. Ut ut omnis.", "Rem ut autem sint ratione magni quos. Omnis voluptatem suscipit earum debitis corrupti. Eligendi aliquam voluptas et rem. Corrupti magnam fugit.", "Qui molestiae laborum in perferendis dolor eum. Quae consequuntur rerum laborum illo. Voluptatem suscipit accusantium asperiores dignissimos.", "At a molestias dignissimos voluptatem est. Odit odio vitae consequatur totam dignissimos aut nam. Et exercitationem voluptas labore velit. Aut omnis incidunt vero et quo."]