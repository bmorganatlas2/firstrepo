["Enim velit tempore labore eum assumenda. Dolor est modi nostrum non omnis quos. Laudantium atque provident sint. Dolorem ut asperiores accusantium.", "Voluptatem est quo quaerat et ut. Quia officiis tempore sed praesentium similique. Explicabo perspiciatis est atque. Deleniti molestiae architecto.", "Quis est sunt. Sunt nulla repellendus placeat consequatur. Architecto corporis commodi ipsum id voluptatum. Animi earum facilis. Libero quis et officiis aut facilis vel.", "At error vel. Sit quis autem quasi doloremque architecto vitae voluptate. Ut et qui.", "Sed dolor alias porro. Eum odit qui esse corporis. Architecto aperiam sit voluptatum nesciunt quia aut.", "Numquam excepturi eos illo qui. Veniam facere eius mollitia et. Qui cupiditate sunt voluptates praesentium.", "At et deserunt non ipsum. Blanditiis qui rem autem. Sed voluptas eos dicta reprehenderit nostrum sed recusandae.", "Rerum quibusdam cumque. Sunt eaque rerum vitae pariatur explicabo asperiores inventore. Necessitatibus impedit neque modi cupiditate magni. Nisi delectus facilis ipsam nulla.", "Aut qui laboriosam non. Reprehenderit labore est. Et dolor voluptates corrupti. Maiores occaecati nihil."]