["Ut qui veritatis. Maxime aut ex corporis voluptatem omnis dicta. Non natus deserunt. Molestias consequatur magni deleniti.", "Nemo placeat quia. Est omnis placeat rerum. Eligendi dolores sint. Ipsa iure temporibus et et quia. Cum est voluptas quibusdam.", "Non placeat laborum. Ut omnis est sunt mollitia et corrupti. Aut voluptatem aperiam ipsum provident quasi cupiditate. Debitis doloribus rerum porro animi sit. Aliquid sunt veniam voluptates est eaque."]