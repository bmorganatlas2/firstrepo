["Ex harum at. Eaque blanditiis vel in. Dolores corporis maiores voluptatem adipisci velit.", "Animi pariatur sit molestiae ut voluptatem quia omnis. Itaque at sed asperiores. Sit porro officiis dolor."]