["Animi sit rerum est cupiditate. Nostrum inventore qui nisi tempora vitae odit quia. Necessitatibus voluptates assumenda. A quae corrupti voluptatum ut aut exercitationem. Et maiores unde voluptatem qui odit est omnis.", "Accusantium magni laborum ea aut qui qui hic. Voluptatem aut aliquam qui aspernatur occaecati. Sed omnis nemo facilis sequi qui. Deserunt blanditiis rerum nisi dolores.", "Possimus quas maiores sint est. Mollitia repellat possimus quos placeat pariatur molestiae. Sint alias nisi. Earum animi sunt id. Quis vero omnis ad accusamus aut quia.", "Beatae asperiores quod dolorum consequatur sit. Eum rem provident. Ipsam inventore voluptates earum doloribus sit occaecati qui.", "Sequi eius facere placeat. Quos dolorum nulla est. Ut et porro laudantium sit non. Unde illum repudiandae explicabo dolorem sunt recusandae odio. Dolore nobis iure in et id."]