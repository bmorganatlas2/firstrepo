["Non rerum magni. Laudantium sapiente tempore. Quaerat consectetur doloremque. Nobis qui dolorem perspiciatis vel magnam. Consequatur explicabo veniam perspiciatis.", "Ea consequatur fugit cupiditate saepe quisquam magnam iste. Architecto soluta est sunt labore impedit in. Quaerat ut ab ut enim autem.", "Hic nihil laboriosam adipisci exercitationem velit omnis. Dolore id numquam tempora. Et corrupti illum eum qui eligendi doloribus velit. Assumenda dolores architecto autem atque corrupti qui voluptate. Laborum id distinctio.", "Voluptatem aut culpa blanditiis voluptas enim alias explicabo. Nulla ullam voluptatem ipsam. Mollitia qui eveniet consectetur placeat quae aut. Possimus hic voluptatum voluptas. Ducimus tenetur culpa.", "Sunt explicabo rerum facere iste. Ratione ut dolore. Aut sit commodi id aut. Eius laudantium quo iusto velit non magnam.", "Dolorem magni earum vitae temporibus non est. Sapiente suscipit eligendi aut ut neque quos. Deleniti eos voluptatem. Necessitatibus qui beatae perspiciatis inventore omnis incidunt voluptatem.", "Itaque culpa est. Et iusto ut quas recusandae laudantium commodi consequatur. Quaerat assumenda impedit eos et necessitatibus ea.", "Accusamus qui corrupti aut aliquid doloribus. Non itaque quaerat corrupti quidem. Rem amet laboriosam."]