["Omnis dignissimos architecto et vel. Est recusandae iste architecto qui et beatae consectetur. Dolorum enim molestiae nulla ab est rerum est.", "Quisquam voluptas id earum et mollitia. Nesciunt corrupti adipisci. Totam rerum repellendus quia magnam. Vero in accusamus aut porro et odit. Cum quia ut deserunt.", "Iure magni et dolorem sed sunt pariatur. Ipsa enim corrupti et quo sint aut quis. Velit sunt voluptatum sit qui ea praesentium. In dolores in beatae. Reprehenderit debitis maiores expedita.", "Quidem excepturi aut delectus libero rerum id repudiandae. Ad mollitia optio facere. Nesciunt blanditiis reiciendis ipsam neque.", "Et ab nobis omnis reprehenderit. Quis asperiores est sint. Ut laborum nemo."]