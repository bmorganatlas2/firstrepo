["Natus et quis aspernatur non tempora sunt veniam. Iste quam accusamus omnis quos id aliquid dolorum. Accusamus quia ad hic cum.", "Qui est voluptas placeat aut voluptatem aut aut. A nulla vel. Iure quo voluptates velit et laboriosam omnis quis.", "Laborum quod nesciunt suscipit. Nihil ut id consequuntur perspiciatis ab voluptate. Non et qui eum a non debitis.", "Velit voluptatem similique sed quisquam. Quia animi repellat maiores asperiores dolor. Qui temporibus excepturi est voluptates nihil. Mollitia assumenda aut veniam aut voluptatem omnis. Eos voluptate earum laborum ipsam.", "Quibusdam molestiae dicta aspernatur doloremque vero non blanditiis. Illum sunt perspiciatis sapiente. Illum eaque a iure omnis. Dicta dolor et qui aliquam. Beatae iusto possimus.", "Suscipit eos deserunt at. Similique dolorem nemo perspiciatis aliquam hic. Quidem ab maxime perspiciatis. Commodi velit dignissimos quo unde. Quod eveniet quos omnis et.", "Qui quia et magnam aut atque nostrum facilis. Occaecati libero cupiditate. Et tenetur sunt consequatur ut eum enim excepturi.", "Vitae reprehenderit voluptatem dicta quidem et veniam. Ratione soluta voluptas commodi non atque nobis fugiat. Rerum delectus nisi ea voluptas omnis necessitatibus.", "Provident reprehenderit ad. Molestiae temporibus dicta suscipit eos culpa. Minus sit ducimus ipsam dolorem quia nihil. Quod temporibus cupiditate quas ea veniam est rerum. Consequatur suscipit delectus nulla et labore."]