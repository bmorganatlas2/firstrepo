["Dolor veniam et necessitatibus modi laboriosam rerum quo. Ab nulla in soluta quia est eaque doloribus. Et cum labore tempore. Voluptatibus consequuntur ab distinctio.", "Optio error nesciunt et vel. Velit iste qui deleniti sint aliquid quibusdam. Et accusamus itaque et laborum corrupti. Quod perferendis laboriosam aut est veritatis deserunt quas.", "Molestiae doloribus in qui perspiciatis minima natus non. Dolorem non omnis. Dolorem qui mollitia consectetur. Assumenda laudantium alias.", "Accusamus ipsa non voluptatem aut suscipit. Eligendi voluptatum consequuntur numquam quia nesciunt omnis sunt. Deleniti sed perspiciatis aliquid illo incidunt laborum.", "Quae earum tempora nostrum dolorem beatae et autem. Incidunt reprehenderit aut nihil porro et. Consequatur et quasi.", "Magni earum minima expedita repellendus praesentium odio nobis. Quas sed ipsam eum est. Aut eveniet ut architecto quo magnam qui molestiae. Sint consectetur veniam quam sed praesentium iure.", "Repellat minima aspernatur aliquid. Voluptatum iste et voluptatem porro odio omnis provident. Debitis minima fugit. Voluptate repudiandae eius voluptas.", "Repudiandae velit id autem omnis. Eum quia consequatur. Est eaque et repellendus vero."]