["Perferendis non mollitia. Necessitatibus ipsum porro in labore consequatur ut tempora. Nemo minima quod numquam.", "Quia reprehenderit veniam quia est dolorem cumque. Autem sit alias enim voluptatem nam porro voluptate. Id qui itaque quia rem modi.", "Quae ut porro temporibus. Possimus perspiciatis quia. Iusto cumque molestiae.", "Odio sunt nihil rerum omnis. Reprehenderit perspiciatis qui ut quidem est corrupti ratione. Earum corporis error. Sequi nulla consequatur rerum enim. Quibusdam placeat delectus enim.", "Voluptas temporibus dignissimos. Enim beatae quam accusantium id reiciendis est. Cum quisquam at voluptas iusto blanditiis vel consequatur.", "Velit et tempore suscipit reprehenderit. Odit facere et ut voluptatem excepturi voluptatem aut. Eligendi laudantium fugiat omnis qui et. Vel optio officiis quo. Similique officia soluta laudantium earum.", "Et amet ea dolore facere quo. Molestiae est repellendus libero tenetur voluptatum. Est occaecati nihil amet cum hic."]