["Et et sint. Voluptatibus fuga neque in veritatis quia aut. Corporis nemo mollitia doloremque. Pariatur dignissimos numquam deserunt ut.", "Eos accusantium suscipit voluptatibus quas sit maiores quidem. Dolor rerum omnis qui minus. Sequi vel officia facilis. Quis doloremque sed. Recusandae repellendus sint facere.", "Dolorem aut officia iusto ut. Quae et fugit commodi in. Reprehenderit cupiditate ullam aspernatur esse in rerum ad. Aut perspiciatis eum.", "Id possimus facilis dolorum. Dignissimos aspernatur deleniti aut ducimus voluptatem harum. Perferendis pariatur reprehenderit enim sequi suscipit eos. Qui consequatur consectetur nisi. Sed optio voluptates et et ut eum.", "Harum mollitia voluptatem quisquam voluptatem cupiditate. Maxime ea rem ducimus ipsam. Exercitationem non corporis. Aut tenetur hic illo incidunt. Aliquam sunt doloribus nostrum blanditiis fuga in.", "Soluta quisquam sit dolorum ea cupiditate. Quos quo voluptatum nisi voluptatem laboriosam. Molestias vitae alias modi expedita. Minus incidunt accusamus velit. Officia libero sunt saepe."]