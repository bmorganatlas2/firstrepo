["Dolorem nihil et autem quod perspiciatis qui itaque. Esse nulla dolores quas id dolorem optio et. Id harum ab velit aperiam expedita molestias. Libero aut dolores. Quisquam placeat et qui facilis vitae ea officiis.", "Velit deserunt commodi et eum tempore tempora fugit. Mollitia possimus occaecati commodi alias impedit tempora consequuntur. Repellendus facilis voluptas perspiciatis sed.", "Pariatur eos incidunt. Magni culpa ea maiores. Fuga explicabo consequatur accusantium nemo quia quis qui. Voluptates ducimus doloribus aut.", "Excepturi exercitationem praesentium quis molestias totam. Commodi enim quam voluptatibus quaerat. Veniam est molestiae iusto itaque ut ut repellendus. Non tenetur enim dolore voluptatibus. Omnis sequi iure.", "Cupiditate omnis recusandae dolorem ducimus. Voluptates nobis labore est. Tempore sit sequi unde nobis. Voluptatem veniam ratione qui soluta enim voluptates a. Nobis esse sunt.", "Dolor a nam. Voluptatem at velit sit accusantium aperiam cumque. Sit ea in atque nostrum ad minus et.", "Ab ipsam delectus eum. Sunt sapiente ipsum ratione eaque enim tempore. Cupiditate totam autem quam nihil. Rerum optio rerum et blanditiis eos voluptatem. Maxime nulla magni excepturi facere cupiditate.", "Odio ducimus iure amet et voluptatem aspernatur. Aut incidunt id perferendis. Distinctio eos a omnis quisquam non vel. Consequatur repellendus dolorem harum ex exercitationem cumque qui. Vero minima numquam excepturi.", "Expedita nostrum est sequi doloribus dolores. Occaecati voluptatem consequuntur molestiae. Voluptates cupiditate consectetur ex et laborum autem."]