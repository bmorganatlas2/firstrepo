["Aut in doloremque non corrupti quis non. Quas ducimus vero iste et voluptas est molestias. Itaque quis quam.", "Nemo quia dolorum blanditiis et tempora deleniti. Quo sapiente est. Nihil molestiae illo eum. Tempore esse eum ut quia sed ullam.", "Autem voluptates eaque perferendis inventore dolorum ipsam ipsa. Cupiditate ad odio tempora aliquid dolores nihil consequatur. Et hic saepe. Molestiae autem vero omnis rem quis at.", "Officiis quo est illum et qui. In sed ea. Assumenda dolor dolorem nesciunt. Reiciendis facere et soluta quia dolorem est eum. Repellat aut est qui velit et.", "Et sunt quos qui molestiae. Praesentium autem enim excepturi accusamus et. Voluptas officiis corrupti incidunt. Eum libero sunt perferendis alias ut."]