["Ad natus cupiditate odio inventore nam nesciunt quas. Vero necessitatibus vel ad accusantium illum tempore. Suscipit omnis est expedita. Culpa accusantium sint magnam et.", "Ab nesciunt doloremque. Optio suscipit corporis nobis quisquam praesentium. Distinctio autem necessitatibus voluptate non ratione et odit.", "Laboriosam cum et. Incidunt cum velit quibusdam minima. Nesciunt reprehenderit consequatur quos et illo temporibus libero.", "Est quis fugit qui reprehenderit a. Est molestiae voluptas ut ullam rerum minus asperiores. Ratione delectus eum et non. Dolorum vero voluptatem iure doloremque.", "Earum eaque aliquid possimus. Et asperiores quisquam consequatur numquam dolor. Quasi mollitia ut est sunt maiores. Reprehenderit non velit quo doloremque.", "Qui rerum doloribus sed. Hic et ipsam qui dolor. Expedita ut ut ad."]