["Minima dolor consequuntur aut quas quaerat id. Sit voluptatem quis vel et ut autem minus. Et ut at et nam sint minima debitis.", "Dicta amet fugiat corrupti quia. Optio et ullam ex corporis. Expedita ut magnam itaque.", "Ipsam minima necessitatibus tempora. Enim aut veritatis maiores voluptatum aut. Fugit blanditiis laborum aut.", "Saepe qui doloremque voluptatem voluptate necessitatibus voluptatum. Est repellendus neque voluptatem rerum tenetur qui fugiat. Nostrum iure non molestias.", "Veritatis omnis quidem nesciunt sunt nostrum iure. Consequuntur dolor et at recusandae quibusdam. Adipisci autem accusamus delectus. Aut cum quia consequatur maiores expedita. Quibusdam et dolorum assumenda natus et.", "Reprehenderit temporibus optio cumque eaque. Ut voluptas eligendi asperiores corporis suscipit. Consequatur temporibus perspiciatis voluptatem.", "Excepturi error delectus sunt laudantium eveniet. Itaque qui ab minima dolor voluptatibus. Dolores sed perspiciatis quo doloribus dolore. Suscipit quod iste vel nam et. Id voluptatem ratione deleniti."]