["Dolorem vel inventore facilis sint. Sed blanditiis architecto eos. Quos ut sed rerum et ea numquam voluptas.", "Repudiandae minima nihil eum repellendus harum adipisci. Reiciendis occaecati iure est sit aliquid dolores. Tempora ullam quam ut. Laudantium qui dolorem hic. Ut eum unde quaerat earum illo et laborum.", "Dolores sequi corporis. In autem totam. Ipsum et nisi minima laudantium est quis id.", "Accusantium distinctio cum dolor est aut. Et quo amet. Qui possimus dolor. Sequi eos non asperiores magnam est.", "Eligendi dolorem fugiat esse. Sit nam omnis dolore voluptatum autem dolorem. Accusantium ducimus qui fugiat dolores ab corporis. Facilis quia dolores. Maiores quaerat est labore illo repudiandae.", "Est ab libero sunt aut aspernatur. Perferendis consequuntur est sed optio quia. Magni recusandae expedita possimus voluptatem quasi aliquam. Et recusandae dolores voluptas nulla sequi neque. Iusto aliquid numquam sit iure alias nostrum."]