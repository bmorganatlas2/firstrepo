["Et debitis autem provident recusandae qui voluptatem. Corporis fugiat non autem commodi labore eos. Ut dolorum qui placeat. Suscipit in voluptas perspiciatis hic qui.", "Facere quam deserunt totam. Numquam minus est. Blanditiis quam velit magnam. Harum laborum eaque maxime veniam reprehenderit aut.", "Quia sint temporibus incidunt dignissimos qui laboriosam corrupti. Aliquid deleniti est animi. Voluptatum a facere. Repellat perspiciatis itaque et laborum ratione. Aut maxime optio incidunt.", "Repudiandae enim et et incidunt sint deleniti. Sunt ut qui et voluptatum. Fuga rerum et aut qui.", "Dolor sunt molestiae beatae consequatur. Architecto expedita est ducimus. Consectetur minus accusamus quisquam veniam quam modi. Exercitationem eum a maiores quo velit est et. Quo nemo soluta illum consequatur."]