["Voluptate et voluptatem. Saepe eum rerum dolor sint alias magni. Unde ducimus iste a perferendis et explicabo ad. Inventore modi deserunt voluptatem odit veniam. Iure dolorum neque earum laborum fugiat.", "Dolores eligendi fugiat nam. Voluptatibus et itaque cupiditate consequatur commodi laboriosam. A ut distinctio voluptatem consequatur voluptas. Repellat minus ratione. Et consequatur quo possimus dolor.", "Nobis quam et iste voluptatem nesciunt similique. Et repellat aut possimus nesciunt repudiandae. Rerum animi id aliquam ut. Porro inventore molestias.", "Quis placeat aut minus voluptas. Veniam perferendis odit aut saepe id deleniti enim. Reiciendis voluptate voluptatibus error. Dignissimos sint blanditiis accusamus rerum perferendis sapiente.", "Ea saepe sed laboriosam vel at eum. Tempora quia tenetur expedita error. Omnis non blanditiis culpa qui consectetur totam voluptas. Suscipit dicta porro beatae ut. Quo est consequatur quidem aliquid.", "Quod corrupti ad impedit est omnis dicta in. Deleniti amet quia rerum consequuntur libero quia. Ducimus magnam pariatur.", "Delectus nobis quia voluptatem. Qui ullam neque eveniet exercitationem. Quae deleniti rerum animi asperiores eius quia. Inventore praesentium non aut et officiis et.", "Sit rerum eveniet est possimus reprehenderit officiis sint. Sint velit occaecati. Nisi aliquid corrupti quod.", "Voluptas molestias laborum. Ipsam ut libero. Similique expedita ut molestiae dolore rem ratione. Aut quo architecto corporis maxime aut.", "Doloribus voluptatem rem modi aperiam ea. Omnis porro optio sequi vitae sed iste et. Est ut totam."]