["Aut quam rem. Officiis dolorem debitis. Sint nisi repudiandae. Maxime eum asperiores velit laboriosam. Rerum quod quia praesentium velit velit."]