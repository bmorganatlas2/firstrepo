["Nulla veniam sed. Recusandae assumenda fugit natus. Amet molestiae hic aspernatur labore commodi unde libero. Rerum aut perferendis laboriosam repellat. In omnis ut pariatur eius qui itaque porro.", "Rerum quia quo magnam. Doloremque impedit nam quos autem. Qui aut et harum modi voluptatem dolor. Odit omnis corrupti rerum. Et inventore qui consequatur."]