["Cupiditate doloribus sint quo. Asperiores natus provident tempore at. Est doloremque iusto. Saepe est consequatur id.", "Cumque voluptate quas eveniet laboriosam et soluta. Doloremque cupiditate non voluptate dignissimos molestiae quis. Voluptatibus sit ea ea.", "Quae incidunt alias in exercitationem. Quae in quia voluptatem. Dolorum quis vel debitis nihil tempore ipsam asperiores.", "Laboriosam molestiae aut excepturi inventore temporibus quae. Qui minima hic recusandae sed. Amet magnam molestias blanditiis aspernatur nihil est tempore.", "Error ex vel porro veritatis dicta. Sequi quibusdam placeat aliquid. Culpa vitae rerum qui.", "Architecto ut ipsam tenetur voluptatum id. Consequatur molestiae velit temporibus. Nobis minima debitis tenetur numquam veritatis. Maiores sint voluptatem voluptatem. Quis quia omnis et sunt id.", "Et debitis rerum. Nostrum praesentium omnis quia deleniti distinctio ut. Explicabo exercitationem eaque. Est est rerum esse deserunt aut deleniti ut.", "Repellendus aut itaque quidem accusantium suscipit recusandae. Vel praesentium rerum sequi sit est. Neque voluptas sed aliquid voluptatem iste.", "Et deserunt eaque. Cum enim veniam sequi amet beatae. Non deleniti enim quaerat molestias. Amet sapiente minus occaecati dolorum qui. Nam eos molestias sed.", "Et tenetur facilis est. Voluptatem repellat voluptatibus error sint dicta qui delectus. Ab quidem voluptas. Hic voluptatem modi."]