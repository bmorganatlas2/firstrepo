["Repudiandae ipsum accusantium animi ut earum. Reiciendis voluptate eligendi labore. Praesentium sit sequi optio culpa. Et illum consequuntur sit. Quis eos rerum et.", "Doloribus earum praesentium quia. At unde pariatur. Nulla fuga nemo enim modi aut illum. In impedit id et. Rerum ut sint id molestias harum a sed.", "Eos suscipit est quia est. Eveniet ratione neque sed. Voluptas exercitationem dignissimos dolor neque consequatur.", "Et deserunt itaque ad earum et. Doloremque tempora non voluptatem quisquam iusto occaecati. Aut iusto voluptas unde quaerat saepe. Veritatis qui ducimus dolor. Eligendi fuga optio nostrum incidunt commodi.", "Sed est sint nulla rerum non. Odio ratione molestiae veniam rerum. Ex ullam aliquam rerum unde dignissimos. Excepturi nam reprehenderit eum esse ipsum. Maiores vitae quas repudiandae non laudantium qui alias.", "Libero velit neque illum aut eveniet. Reiciendis ratione quas dolore eum dolor eos. Voluptas veritatis illum rerum voluptas.", "Harum maiores culpa quia dolor. Tempore numquam magni. Consequatur placeat iure voluptatem voluptates quia. Nisi consequatur non ea suscipit quia non.", "Autem in reprehenderit sapiente cumque doloribus et veritatis. Sed quaerat eius. Nam veritatis quis soluta atque est adipisci. Dolores sed molestias beatae autem sit.", "Corporis tempore atque blanditiis est omnis in. Voluptates voluptatem beatae enim sed consequatur et magni. Amet in dicta atque. Et est quisquam. Deserunt vero dolores ab corrupti illo sit impedit.", "Corrupti harum qui illo natus eos. Nihil harum quaerat autem qui. Et ut repellat sed qui ut autem. Dolore eligendi iure. Est ut veritatis tempore recusandae amet nihil ut."]