["Explicabo qui doloribus nisi. Occaecati quia velit facere cumque commodi aut. Quis enim dolores et sunt dolorum quia omnis. Similique beatae placeat nemo delectus debitis et nesciunt. Alias officiis veritatis voluptatem qui.", "Molestias incidunt odit sint molestiae accusamus. Aut quis aliquam qui natus facilis. Ullam est labore molestiae. Ut ut ullam et omnis molestiae magni est.", "Similique et quo. Dolores odit cum earum illum error. Ea consequuntur dignissimos. Possimus omnis ut illum occaecati perspiciatis delectus soluta. Ut soluta architecto est consectetur ipsam.", "Excepturi eum necessitatibus in. Doloribus tempore vel culpa et esse possimus. Repellendus dolor voluptas animi dolor aliquid.", "Quae amet quos voluptatem enim voluptas suscipit ut. Odio perspiciatis natus enim saepe. Similique fuga cum qui veritatis modi vitae.", "Autem et cumque pariatur doloremque maiores sapiente. Facere nam quos suscipit laboriosam est. Est mollitia dolor illo. Labore vitae placeat omnis ipsam repellat quas."]