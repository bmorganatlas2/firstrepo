["Odit quibusdam ad enim nihil explicabo. Consequatur dolor repellat voluptatem. Laborum consectetur nulla consequuntur. Consequatur reprehenderit sit sed.", "Officiis quis vel sint aliquid dicta est. Facere aut labore sint omnis excepturi amet nisi. Itaque quae quidem iusto maxime. Eius maxime qui sed nihil id vitae. Ipsam maiores non placeat sequi voluptatem consectetur.", "Enim animi quaerat a aliquam tenetur magnam explicabo. Et blanditiis aut velit. Aut suscipit ut velit sunt eos ut id.", "Culpa est quo porro. Rerum molestiae beatae assumenda iste ipsum. Vitae id ipsam et ut quia qui.", "Fugiat neque voluptates voluptatem. Et non consequatur quisquam ipsum debitis sequi. Exercitationem eligendi nesciunt possimus aliquam et. Alias asperiores minus facere quaerat consequatur est.", "Natus rem quo. Eligendi fuga dolorem. Reprehenderit illum non voluptates aperiam adipisci.", "Eaque id iusto sit sed aspernatur nihil provident. Fugit ut nulla quis. Velit aut sint aut nihil tempora voluptate. Ducimus voluptatum inventore. Asperiores eos quis aliquid eveniet.", "Libero sed suscipit et porro ut eum. Temporibus veritatis similique. Neque reiciendis qui accusamus tempora aut quia perferendis. Consequuntur qui animi dolores quos cumque omnis.", "Et deserunt quam corporis reiciendis repudiandae quas quidem. Ut sapiente velit ea voluptatibus suscipit. Saepe expedita consequatur."]