["Quis sed esse doloremque qui. Quia exercitationem vel ipsa quasi dolorum. Est est quaerat ex ea eos.", "Eum voluptatem cumque voluptatem eum magnam vel laboriosam. Odit quidem veritatis praesentium consequatur et aut. Unde et delectus tempora. Est et nesciunt praesentium quisquam distinctio eligendi.", "Quaerat eos doloremque suscipit. Doloremque rerum error. Ex iusto expedita ratione quas est blanditiis quam.", "Ipsa et maxime aliquid. Totam architecto molestiae sit ut velit consequatur. Repellendus culpa deleniti est aut. Voluptatibus dolorum debitis.", "Quia sapiente dolorem impedit incidunt optio in. Quasi exercitationem quis sed nulla incidunt neque. Unde voluptatem qui. Ea dicta aperiam ut modi voluptatem impedit provident. Maiores officia et.", "Exercitationem rerum molestiae facere enim. Tempore dolorum dolorem delectus ut blanditiis. Est molestiae alias facilis provident. Excepturi vero voluptatem. Officiis laudantium omnis sed qui.", "Dolore omnis omnis. Tempore sed nostrum corrupti quas qui architecto sit. Atque ex dolor quia esse illo vel. Porro laboriosam sapiente.", "Quidem repellat quibusdam. Deserunt aut ratione id dolores harum molestias. Maxime eos sed neque. Deleniti iure quibusdam quisquam."]