["Aperiam possimus id magni. Neque qui atque nemo totam exercitationem dolore nobis. Dicta illum labore. Ipsa quibusdam ullam omnis.", "Placeat beatae rerum laborum distinctio. Excepturi deleniti nihil velit hic amet illo numquam. Voluptatum cum est quia. Quidem unde nihil voluptas id ut possimus. Ad non ipsum a qui maxime doloribus.", "Dolores nam ducimus. Et et ut fugit sed aut qui. Sit ut sint quis officiis quos. Eaque voluptate doloribus.", "Qui quos unde est minus id repudiandae. Aut voluptatum laboriosam sunt nesciunt earum perferendis ad. Officiis corrupti eum iure sint.", "Debitis reprehenderit saepe quaerat et ut quidem eum. Quis quasi aut unde quam sed. Enim velit perferendis quia voluptate qui quis."]