["Sequi alias voluptas voluptas vel blanditiis corrupti pariatur. Porro ducimus reiciendis cupiditate. Quia sint minima ipsam. Non quasi rerum.", "Itaque cumque tempora. Qui officiis adipisci fugiat commodi consequatur quibusdam. Iure vero voluptate nihil accusamus at consequatur.", "Sit itaque est optio repellendus eos. Blanditiis voluptas ut praesentium nemo et quis. Aspernatur et voluptatem veritatis nam quod. Officia sapiente architecto eaque ut quia eos enim. Culpa sit voluptatem."]