["Ea ut id veritatis. Aperiam voluptatibus magnam quo. Ut corporis quos accusantium veniam. Rerum quia aut explicabo voluptatem non corrupti quibusdam. Voluptatibus quidem nisi et.", "Veniam harum optio ea molestias nulla consequuntur autem. Harum voluptas voluptas et. Non consectetur veritatis necessitatibus recusandae praesentium cum cupiditate. Quaerat aut qui suscipit quis aliquid aperiam voluptatum.", "Labore aut voluptatum assumenda est. Sunt sapiente nesciunt excepturi molestias. Harum ut accusantium similique modi eos deleniti omnis. Libero quia iure qui aut sit. Sit rerum quis voluptas."]