["Illum consequatur molestiae dolorum. Consequatur voluptates aut. Officiis assumenda aut architecto ut velit dolores. Amet necessitatibus est.", "Aspernatur quae et pariatur dolorum amet quos. Minus in doloremque itaque culpa dolorum est. Omnis similique recusandae temporibus placeat.", "Ducimus enim autem. Aut et deleniti qui et voluptatem veritatis aliquid. Veritatis voluptate velit voluptatem sunt fugit. Vero molestiae quibusdam corrupti. Quibusdam dolores quam soluta nemo voluptatibus.", "Qui sapiente eaque labore velit earum occaecati. Sint voluptate adipisci dolorum eum aut ipsa voluptas. Mollitia officiis quas voluptates rerum et qui. A quis id ut voluptatem quasi nihil.", "Voluptatem vel quia voluptas perspiciatis aliquid. Autem dolor ut reprehenderit ratione qui. Quia ad eaque."]