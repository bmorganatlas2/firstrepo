["Amet consequatur dolorem nobis est. Ad sunt fuga. Voluptatem voluptatem esse voluptas quia facere vitae. Rerum consequatur non non quis."]