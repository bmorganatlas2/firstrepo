["Numquam dolorum hic eos non. Sit non voluptatibus. Dolor quisquam repellat odio et.", "Magni in assumenda. Quo tenetur est quas. Adipisci consequatur amet sapiente reiciendis. Voluptatum porro laboriosam magnam sed.", "Aspernatur rem dolores. Iste illo error. Voluptatibus tempora exercitationem quas dolores atque dolorum sed. Cum nihil accusantium.", "Voluptate consequuntur est. Dolorem voluptatibus placeat excepturi architecto est magni. Eius deserunt in iste perferendis sint aut aut. Velit qui est id natus.", "Soluta id commodi dolorem eius ut sit. Rerum molestias ea. Eius corporis quia eum molestias impedit qui. Atque sapiente est cumque sit rerum. Et animi veniam.", "Harum rem voluptas dolores dolore voluptatem. Nesciunt similique iste. Nihil reiciendis deserunt autem est eos dignissimos quis.", "Optio ea esse omnis. Excepturi maiores consequatur natus ipsum aut. Non quis reiciendis est aliquam doloribus et.", "Odio et sit voluptatum autem officiis quia. Saepe natus corporis porro ullam quibusdam. Ducimus beatae ut earum quisquam omnis et.", "Numquam distinctio ut doloremque eius quia placeat. Eius voluptatibus placeat error. Eos odio corporis ipsa. Quia eos magnam in. Doloremque animi molestiae ad."]