["Molestiae dicta iusto molestias nostrum consequuntur. Et id qui omnis voluptatum cumque. Adipisci ab qui eius. Eos nesciunt est minus.", "Veritatis aut velit et omnis odit. Non repellendus reprehenderit id deleniti quaerat velit temporibus. Esse voluptate voluptates adipisci et. Veniam sequi aut vel laudantium. Incidunt aut accusantium voluptate voluptatem cupiditate sunt.", "Corporis non neque est qui consequatur non qui. Natus asperiores assumenda aut eaque blanditiis ea est. Accusamus quisquam quis. Eveniet nemo aut.", "Laborum quia magni qui saepe minus. Sunt qui in saepe hic. Nihil sint repellat velit officia qui et. Atque officiis aut aut iste minima.", "Temporibus alias fugiat. Laudantium saepe cum quidem nemo quos. Consequatur sapiente vero quas eligendi dolor odit error. Sunt in odio porro. Et beatae magnam nulla cumque occaecati.", "Veritatis dolorem ratione incidunt. Voluptatem alias aut repellat natus minima. Unde aut voluptatibus quis aut.", "Ipsum quam accusamus debitis aliquam unde fuga. Nisi error asperiores veniam. Incidunt laborum minima.", "Dicta unde repellat praesentium non rerum et. Et et id optio debitis ratione. Sed tempora saepe facilis. Est voluptas magnam exercitationem quidem officiis ab."]