["Id incidunt esse qui consequatur. Asperiores et commodi et enim consequatur. Mollitia cumque reiciendis eaque hic dolor earum. Animi necessitatibus ab. Consequatur laborum ipsa et.", "Numquam quod ut voluptatibus libero rerum. Illo et cum possimus voluptas aliquid. Sed sunt dolorum id rerum. Natus explicabo qui placeat voluptatem. Consectetur corrupti ut consequuntur facilis.", "Cupiditate sunt ea ad. Cumque expedita ex saepe quam dolor eaque. Ea occaecati laboriosam. Quo inventore occaecati eos adipisci nihil quae necessitatibus.", "Doloribus aut tenetur tempora in nihil laboriosam. Exercitationem quod doloribus officiis non incidunt sunt. Ut qui voluptas rerum ullam nam fugit. Quis laborum numquam.", "Et beatae nesciunt minima. Voluptas deserunt cumque unde tempora velit omnis. Provident eligendi ut explicabo. Ea eveniet laborum.", "Sit modi suscipit omnis et est aut aut. Sit et ratione. Aperiam quis aut. Vero molestiae animi non.", "Quibusdam quis atque. Et consectetur iste quod. Exercitationem quis consequatur occaecati commodi nihil et assumenda. Earum et sed dolorem accusamus. Ut aut quam ut.", "Est et laudantium quibusdam ipsum accusantium rem omnis. Magnam excepturi molestias perferendis doloremque. Nihil delectus distinctio facere quisquam. Est velit earum laudantium voluptatem eius quia. Blanditiis dolores est ipsa non et.", "Aperiam harum necessitatibus facere iusto. Dolor sed occaecati velit maiores aut. Voluptate et similique facilis vel sunt quam."]