["Numquam ut odit deleniti quo. Aliquid illo necessitatibus enim aperiam sit. Enim sint nisi nihil.", "Consequatur molestiae sed aliquam. Sit dignissimos harum ratione doloribus laboriosam quam. Et ea recusandae voluptatem. Maiores tempore ut natus nihil similique.", "Eum quaerat veniam. Quis facere incidunt dolor nam laboriosam porro. Non delectus numquam. Corporis voluptatem quis sed et. Minus veniam est perferendis sint est autem.", "Et cum dolorum est modi. Perferendis nihil porro commodi labore ea. Tempore sed ut cum. Voluptatem est soluta.", "Sit autem amet tempora. Molestias autem totam quod neque qui. Commodi totam molestias illum quaerat nihil id. Dolore accusamus perferendis.", "Adipisci ut voluptas omnis atque totam qui. Ut eligendi quidem corrupti. Eaque natus et ea voluptatibus laudantium veritatis. Magni et sed excepturi fugit id."]