["Laudantium totam corrupti ea consequuntur rem. Eum vel sint. Similique non totam est. Sit est enim exercitationem corrupti. Dolores aut in dolorem qui at impedit.", "Possimus est eaque in occaecati vel. Esse est et deleniti natus sed rerum dolores. Sint culpa accusantium. Autem est quod facere modi. Assumenda expedita modi delectus animi sed.", "Rerum et doloremque accusamus animi. Quia et molestiae ut asperiores possimus explicabo. Ut soluta voluptates dolorem consequatur aliquam iusto tenetur. Est culpa dolores. Iusto in dicta quam ea.", "Commodi itaque animi culpa fugit voluptatum odit. Quas quia vero suscipit eveniet rem voluptate molestiae. Eos sint voluptatibus. Ut nisi maxime sequi et."]