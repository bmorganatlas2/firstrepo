["Placeat dolorem voluptatem. Voluptas reiciendis culpa exercitationem ab. Aut reiciendis aspernatur.", "Eligendi magnam quos itaque ullam. Quis qui dolores molestias et veritatis et qui. Esse sequi aperiam ut rerum eos aut voluptatem. Possimus dolor nesciunt eos quibusdam eum. Et aut libero a earum assumenda doloribus quis.", "Voluptatem vel assumenda eos exercitationem nihil et aut. Voluptatum voluptatibus temporibus quo quisquam fuga. Cupiditate animi nisi et aut enim occaecati rerum. Veritatis nobis quaerat quis quae temporibus amet voluptatibus. Porro laboriosam voluptas culpa ullam sed.", "Reiciendis qui ut voluptatibus. Facilis nihil error in distinctio eligendi. Eaque voluptatem facere voluptatem. Quia aperiam pariatur accusamus magni. Aspernatur veritatis tempora iste sed reiciendis.", "Consectetur in blanditiis ut vel laudantium sapiente omnis. Debitis quis dolore esse. Quam quidem dolorem ipsam."]