["Rerum eum quos id doloribus possimus ipsam. Consectetur fugit ad ab modi. Optio nihil est et id dolor minus ut. Odit vel iusto possimus qui voluptate quod.", "Autem dolorum eaque reprehenderit ut ut. Fugiat quia aut rerum. Totam aut aut ipsum deserunt. Ut et voluptatem. Voluptatibus possimus eius est molestias quae."]