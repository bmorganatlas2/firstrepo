["Quo deserunt ea ducimus enim. Voluptatem consequatur ipsa. Voluptates enim libero ab a. Id modi sint consequatur nam. Aspernatur ea molestias aut dignissimos quaerat.", "Vitae similique dolorem. Velit laboriosam quod aut. Et quibusdam ut et. Praesentium sit sed. Sequi illum voluptas.", "Consequatur tenetur aperiam dolor sapiente qui maiores optio. Temporibus sunt impedit quidem odio amet harum. Eos magnam similique. A accusamus praesentium. Sed quibusdam dolores."]