["Quos voluptatem quisquam. Omnis cumque ipsum sequi aut ut dicta aliquid. Voluptatem ea voluptatibus quam.", "Et omnis recusandae. Totam ea suscipit. Doloremque sit sed ratione eius expedita saepe et.", "Ut voluptatibus non praesentium temporibus reprehenderit qui ipsum. Error delectus enim doloremque. Et iusto perferendis perspiciatis eaque rerum et voluptas."]