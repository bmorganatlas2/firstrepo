["Molestias quia est amet officia voluptas exercitationem. Reiciendis sunt aliquid nostrum magni illo. Praesentium numquam esse ea tenetur aut quasi id. Ratione illum et eaque quia rerum. Nisi accusamus et voluptas.", "Neque sit in suscipit. Quia necessitatibus omnis optio a. Non aut sed mollitia quia et maxime sint.", "Qui maxime et qui ipsa. Deserunt nam nihil. Aut soluta sunt asperiores ratione quibusdam. Expedita qui aliquam aut non repudiandae. Illum sed error quod cupiditate vitae odio."]