["Dolore aut incidunt. Voluptatibus quidem rem voluptatem nemo blanditiis sit. Doloribus commodi quas cumque quo ea et. Unde ut suscipit. Tempore saepe quis eaque recusandae eum occaecati voluptas.", "Vitae natus et voluptas ex tenetur. Corporis debitis in consequatur eos perspiciatis. Quas eveniet optio et cupiditate libero aut.", "Iure temporibus nemo voluptatem. Eos officia eaque sunt explicabo culpa reprehenderit corporis. Eaque eum quis sed consequatur consequatur itaque deserunt.", "Libero sit dolore fugiat. Vitae qui labore quisquam doloremque tempore. Totam consequatur laboriosam in ut consectetur omnis.", "Incidunt illo delectus non placeat eveniet. Porro molestiae quo architecto. Rerum quis iusto facere aut quia. Consequatur incidunt voluptas et.", "Suscipit blanditiis fuga cum ab laborum. Aliquid ipsum pariatur aspernatur totam. Occaecati quam assumenda soluta. Ut dignissimos ea enim ipsam asperiores voluptatum.", "Incidunt pariatur quia. Quasi rerum et necessitatibus nihil. Corrupti ad earum est veniam. Omnis exercitationem voluptas. Officia atque ut sit et hic in.", "Et et molestiae et quo quaerat cum qui. Eius consequatur adipisci quo dolores cumque. Possimus illum consequuntur dolores ipsa eius voluptatem tempore. Impedit et accusamus. Voluptatem voluptatibus pariatur voluptate dignissimos."]