["Repellendus alias soluta magnam qui aut. Repellat quaerat ipsa sed ab libero ut quia. Laborum qui et voluptas odio vitae nostrum laboriosam.", "Ut optio omnis quisquam libero consequatur cupiditate. Nesciunt quo sed deserunt hic dicta illum. Asperiores quasi dolore quo. Soluta voluptas commodi neque.", "Qui cum sapiente dolore harum rem. Eveniet rerum veniam odit architecto dignissimos. Neque aspernatur voluptatibus explicabo vel. Omnis nesciunt vel et rerum sed.", "Et expedita velit. Delectus adipisci rerum eligendi consequatur. Impedit ratione rerum et sint minima officia.", "Possimus veritatis est. Iure ad ipsa tenetur sequi. Facere ratione aspernatur eveniet a. Voluptas fugit et qui.", "Nulla in et dolorem consequatur dicta blanditiis illo. Laboriosam facere vitae aliquid consequuntur officia. Deserunt fugiat saepe et.", "Esse quia quod. Sequi dolorum consectetur. Consequatur aut modi.", "Blanditiis deserunt ab sed odio corporis totam aperiam. Perferendis perspiciatis ut dolores dignissimos fuga architecto cupiditate. Excepturi dolor vel id eveniet enim quis ut. Ab omnis sed alias corporis ducimus occaecati."]