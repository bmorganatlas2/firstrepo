["At ab illum sit consectetur expedita rem. Architecto iure et illum quaerat debitis. Commodi maxime praesentium corporis. Magni qui similique neque. Molestiae fuga est tempora numquam voluptatem nulla commodi.", "Necessitatibus facere natus corporis quia doloremque libero rerum. Soluta amet nostrum fugiat perferendis atque aut. Dicta soluta et qui. Aut quod sint nam.", "Quae sunt repellat. Et voluptas autem. Doloribus eos eum assumenda dignissimos suscipit. Eius eveniet est dolores impedit praesentium."]