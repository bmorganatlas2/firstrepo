["Molestias eos ab aut maxime. Occaecati veritatis ut quasi porro praesentium modi voluptatem. Cumque nobis ut.", "Magni in voluptas eligendi sit dolores. Iure ipsum veritatis voluptatem aut molestias sequi. Qui eos earum. Ea quisquam et occaecati.", "Quidem laudantium velit dolorem doloremque. Autem labore qui. Magni reiciendis repellendus."]