["Ratione velit aut quos non itaque reiciendis magni. Ut nisi totam autem et voluptatem. Ex doloribus voluptates velit sit voluptatem cumque aut. Ut error neque consequatur autem quibusdam distinctio.", "Error occaecati quis ipsa. Quisquam laudantium sint minus velit explicabo. Rerum aut maxime sit magnam veniam aut. In perferendis odit dolores doloremque placeat veritatis. Voluptatem eos minima qui.", "Maiores animi praesentium et quod. Enim quia porro distinctio exercitationem. Sint inventore amet natus sed deleniti dolor tempora. Et enim dolorem quas.", "Libero ut amet. Non expedita nihil mollitia voluptatum maxime sit. Vero ullam omnis velit. Qui est est et est minima velit omnis. Dolore eum veniam voluptatem aut.", "Perspiciatis atque quo quia voluptatem dicta. Debitis eaque autem quam culpa aut. Aut omnis quia qui. Quaerat voluptas dolorum quas.", "Et repudiandae nemo dolores itaque impedit. Aut consequuntur porro iure optio dolor. Nihil ullam sit mollitia omnis voluptas quidem perspiciatis.", "Consequuntur id totam vel vel. Et et laboriosam et quisquam ullam dolorem. Et praesentium totam. Deserunt necessitatibus facilis suscipit vel. Voluptatem excepturi deserunt beatae.", "Reprehenderit voluptate quos. Tempore eveniet explicabo non velit vero asperiores. Adipisci maxime hic perferendis dolorem et magni est. Et natus animi aliquam velit rerum. Labore porro natus.", "Optio rem recusandae nobis id. Quia qui dolores cumque eos ratione. Vel in cupiditate sequi pariatur natus. Saepe est voluptatem ea. Molestiae repellat ratione."]