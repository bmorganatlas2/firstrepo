["Ipsam impedit et nobis porro quo. Eos sed iste. Earum debitis voluptatem adipisci exercitationem libero occaecati. Accusantium aut voluptates nihil aliquam.", "Accusantium ut aut magni sint unde porro. Quis iure fugiat mollitia dolores possimus omnis. Ea totam reprehenderit. Eos in nobis esse omnis illum.", "Pariatur sit voluptatem eum. Consequatur occaecati accusamus enim. Aut unde ea fugiat quo voluptas iure officiis. Vel qui aut veritatis. Aliquam accusantium possimus eaque qui in dolor tenetur.", "Esse aut expedita. Et voluptate odit ea sed corrupti. Qui in officiis adipisci. Qui aliquid non commodi nihil adipisci est. Laboriosam dicta autem architecto.", "Iure est cum. Libero voluptatem rerum aut dolorem sint. Aperiam eaque recusandae illo atque. Qui laboriosam odio quo fugiat. Dolor ipsa minima dignissimos qui.", "Omnis harum voluptates distinctio. Temporibus odio mollitia voluptas. Aperiam alias voluptatibus et natus. Ullam et est sed quis voluptatibus. Id ipsum eligendi qui quidem nisi.", "Vitae nisi quia. Culpa ab aut reiciendis eum qui officia voluptas. Omnis illo minus ut et fugit sit temporibus. Iure fugit unde molestias nam deserunt excepturi. Quam voluptatem dolores repellat praesentium velit distinctio.", "Ad voluptas nam exercitationem. Doloribus eveniet voluptas. Vero accusamus assumenda harum quibusdam veritatis ipsum et."]