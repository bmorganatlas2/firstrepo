["Nesciunt saepe voluptatem quas cupiditate. Error culpa ut qui. Dolor consequatur nemo culpa voluptatum et sed. Sed et minus praesentium.", "Provident exercitationem ab. Voluptatem voluptatum sunt laboriosam consequuntur aspernatur et. Enim necessitatibus voluptatem. Explicabo culpa aut corporis sunt praesentium."]