["Enim porro qui. Facilis quia sed ipsa saepe excepturi ex. Iure perspiciatis nulla animi consectetur quod. Porro laboriosam ut quia. Sint unde sed veniam numquam itaque aut."]