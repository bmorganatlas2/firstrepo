["Earum officia illum et. Ut est ea. Velit voluptate laboriosam odit numquam quisquam nam consequatur. Facere sed recusandae veniam voluptatem. A esse et sunt temporibus sit deleniti officia.", "Nihil placeat veritatis. Quas sed doloribus maxime. Qui ipsum qui.", "Possimus ex qui. Inventore culpa quia officiis incidunt et. Quia at eveniet qui."]