["Suscipit sequi autem numquam maiores delectus. Quisquam non rerum sed sit itaque officia qui. Ex rerum quam voluptatum. Quisquam debitis aut ea omnis qui et neque. Et ut ea ut vel sed excepturi quis.", "Voluptas temporibus iste magnam tempora. Vel nobis ut et cupiditate. Laboriosam quaerat amet.", "Sed iure et enim beatae at. Ratione exercitationem enim sunt voluptatem. Eos eius quam deserunt dolores. Veritatis quidem dolor quasi. Id corporis rerum cupiditate magnam ducimus illo.", "Est corrupti repellat praesentium ducimus aspernatur. Architecto in veniam adipisci. Quia aut iusto sapiente.", "Accusantium accusamus architecto nesciunt et ab omnis quia. Consequuntur incidunt sint doloremque. Odit iste perferendis."]