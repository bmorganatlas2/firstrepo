["Assumenda vero sequi ea sit dolores enim. Quisquam quia magnam sequi voluptatem qui enim. Error iusto beatae odio. Recusandae non ipsa qui iusto dolorum.", "Debitis quo aut aspernatur alias earum consectetur. Doloribus dignissimos quia beatae tempore quo rem vel. Dignissimos facere nobis illum veniam autem."]