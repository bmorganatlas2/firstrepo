["Qui sint quos. Ipsa rerum quaerat. Eligendi sit iste eaque magnam quod.", "Ut dolorem modi reprehenderit voluptas harum vitae. Officia sint cumque. Sint totam nihil ex tempora consequatur quibusdam harum.", "Iusto consequatur est non voluptas eligendi. Sit et consequuntur adipisci odio. Quam ut est. Quo exercitationem et dolores pariatur officiis."]