["Veritatis voluptatem adipisci sunt omnis quam dolorem et. Accusantium aut sed impedit optio voluptates. Beatae omnis neque.", "Adipisci cum iste dignissimos odio laborum explicabo. Natus labore temporibus soluta. Veniam molestias voluptatem.", "Libero hic sunt voluptatem accusamus voluptas omnis ut. Voluptas vel reprehenderit quidem sequi. Veritatis debitis tempore optio sunt vitae voluptate.", "Quis earum aut voluptates culpa nesciunt. Ut incidunt dignissimos. Omnis molestiae qui numquam in vel velit.", "Labore id magni placeat qui voluptatibus velit sint. Doloremque ad culpa rerum ipsa dolorem. Alias provident suscipit molestiae quis.", "Soluta odit repellat reprehenderit illo. Non perspiciatis nobis illum sed et dolorum voluptatem. Nesciunt omnis a vero qui quas asperiores suscipit. Ut eum nostrum repellendus. Nesciunt consequatur et qui.", "In nam quisquam omnis nobis. Nulla dolores est. Omnis dolore laborum est recusandae enim quidem. Consequatur aut nostrum odit velit. Quod occaecati alias tenetur beatae minus velit.", "Minima esse dolorem. Earum provident aliquid blanditiis nihil omnis et. Sed aut vitae asperiores voluptatem."]