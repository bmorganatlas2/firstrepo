["Non est et. Animi consequuntur laboriosam aut omnis dicta fugiat sed. Error cum est quisquam. Sint odio voluptatem ut sequi. Enim omnis minus itaque numquam nihil rem harum."]