["Dolorem quis id qui autem ab sapiente rerum. Voluptatum ut dolor quis omnis quasi. Sapiente rerum autem dolorum eum quo quod et.", "Quia sed et sed. Quia et qui. Fuga veritatis et sed tempore autem voluptatem."]