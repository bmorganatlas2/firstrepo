["Repudiandae doloremque est modi voluptatem. Beatae repellendus illum facere corporis quasi repudiandae. Nihil qui dolore magnam ratione fugiat illo. Maxime quia quis.", "Totam quo sint eum rerum et velit voluptates. Odio eos quae recusandae veritatis. Quia labore et reiciendis. Voluptatem consequatur nam. Qui dolor in vero sint.", "Sunt dignissimos voluptatibus dolore architecto. Qui quis vitae in sequi error. Error numquam omnis. Molestiae impedit ratione adipisci suscipit illum. Excepturi sunt laborum omnis quod et."]