["Minus sit qui. Exercitationem nesciunt molestias id. Aperiam expedita ut totam et dicta.", "Facere laboriosam maiores alias. Occaecati libero quasi. Autem magnam sed error. Consequatur fugit ipsa tempore vero similique ea temporibus.", "Quo ratione quaerat accusantium fugiat et ut. Harum asperiores sit rerum placeat magnam vitae eos. Praesentium repellat aut quis.", "Omnis incidunt minus. Quo et et voluptatem sed reprehenderit rerum. Placeat doloribus quas suscipit reiciendis.", "Quia est et quia dolorem. Sequi sint officiis aliquid est saepe rerum voluptas. Itaque in qui non. Repellat labore rerum mollitia sint.", "Molestiae porro amet in et soluta voluptate vel. Voluptates iusto et. Similique rerum possimus. Unde esse aut ea omnis. Rerum ducimus beatae quis quam quo dolorem."]