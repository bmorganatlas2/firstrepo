["Id dolorum vitae minus aut. Sequi illum illo et consectetur. Minima consequatur ad cum et. Laudantium pariatur exercitationem nemo nostrum quisquam.", "Cum repudiandae at. Tempore consequatur officiis vel placeat. Exercitationem inventore neque qui itaque nesciunt distinctio. Vel impedit et sed cumque quam exercitationem.", "In quis alias culpa. A voluptas quidem atque. Non soluta laborum quos mollitia nulla cumque aut. Et provident facere accusantium molestiae voluptatem placeat.", "Nihil quis voluptate omnis laborum ipsa. Voluptatem suscipit tempore sit. Aut architecto enim qui quos sapiente esse.", "Dolorum odit expedita nihil. Velit eaque distinctio tenetur animi quia earum. Reprehenderit alias commodi.", "Qui rerum cum incidunt. Assumenda tempora consectetur incidunt dignissimos et nemo necessitatibus. Vel ad autem possimus saepe ut rerum suscipit. Ducimus eveniet ut. Est molestiae voluptate.", "Voluptatem ea corrupti ipsam. Dolor in dignissimos enim aut recusandae aut. Adipisci omnis deserunt cum optio ea aliquid ut. Libero non tempore et distinctio veniam nihil quam."]