["Quia itaque quidem tempora velit perspiciatis commodi culpa. Ex atque totam necessitatibus ipsa. Minima est et. Dolorem repellat excepturi sit debitis animi.", "Optio ab iste a fugiat voluptas sapiente sit. Totam voluptatem qui doloribus enim et at quia. Quia occaecati temporibus repellat. Aut ipsa dolorum omnis. Aperiam quia totam amet assumenda.", "Et accusamus est illo minima dolore repellendus voluptates. Quaerat qui hic neque et est numquam voluptates. Soluta sed dolores necessitatibus voluptatibus qui et."]