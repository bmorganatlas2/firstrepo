["Est natus velit. Nihil molestiae voluptatem consequatur. Deserunt commodi quisquam quae magni.", "Sunt minus iste et beatae perferendis animi. Et minima sunt. Aut dolorum culpa amet iure nesciunt incidunt. Necessitatibus labore sint. Commodi eos atque et dolores.", "Ut alias est provident. Suscipit soluta totam eligendi dicta culpa. Quo ut quidem rerum eum tempore consequatur. Porro id fugiat. Occaecati sit similique mollitia eveniet.", "Laboriosam laborum velit voluptas atque mollitia dolore. Ut sit qui. Molestias quibusdam modi. Culpa et et sint.", "Rerum quam commodi animi quis omnis. Soluta sint nisi ratione ipsa quaerat. Error voluptatem tempora numquam est. Molestiae ducimus facilis ab dolore quaerat non.", "Illo sed minus et a quidem est. Molestias id esse suscipit. Omnis explicabo tempora expedita molestiae distinctio nisi quae.", "Voluptate magni rerum alias aut consequatur libero hic. Qui aut labore eius. Quia aut eaque quos aut consequatur. Doloremque occaecati asperiores est. Praesentium distinctio nihil deserunt quia recusandae cumque commodi.", "Repellendus voluptatem nobis ut et suscipit. Et perspiciatis at quis saepe mollitia architecto. Ipsam quaerat asperiores quisquam quia saepe.", "Quos nesciunt corporis eveniet perspiciatis delectus facere. Veniam asperiores autem placeat aspernatur sunt dolor est. Repudiandae voluptatem incidunt dolores minus earum.", "Quibusdam veritatis voluptas eum qui voluptates ut. Impedit autem alias doloremque. Maxime in et dolorem."]