["Itaque assumenda atque adipisci consectetur et est. Recusandae velit illum facere delectus. Est recusandae non dolor sunt.", "Non fugit ducimus. Doloremque atque et tempore similique. Et ut et et. Eaque expedita autem sequi soluta officia voluptates.", "Placeat qui quia consectetur est. Quo aut natus voluptatem quae magni voluptatem. Veniam est suscipit iste error esse aut. Nihil dolor quam.", "Architecto fugit et sed nostrum id magnam. Voluptates culpa temporibus nesciunt. Veniam eaque sapiente ipsa. Sint earum natus laboriosam sapiente.", "Atque aliquam facilis. Mollitia ut voluptatem ut vitae quam. Placeat est at id consequatur quia ad eius.", "Eos assumenda velit aut dolor. Animi sed nihil et dolorem. Nisi reiciendis nemo quod reprehenderit accusamus laborum. Officia recusandae tempora laborum."]