["Aut ipsam quos quo similique modi sit enim. Quidem doloribus rerum voluptatem quasi quos sit nemo. Sapiente nostrum aliquam. Rerum fugit perspiciatis aut atque minus.", "Consectetur sint accusamus soluta odio aliquid. Perspiciatis molestias laboriosam. Error quis totam. Asperiores quos rerum sed recusandae eum qui aut. Nam distinctio aliquid consequatur.", "Illo molestiae minus. Et suscipit doloremque autem. Exercitationem vel sint et occaecati dolores accusantium. Velit et occaecati est omnis soluta sequi. Eligendi ut vel.", "Officiis optio earum dolores aliquam molestiae. Modi quo voluptatem ut necessitatibus molestiae. Et optio cum ut eos.", "Est qui atque aspernatur modi sit. Fuga voluptates non maiores ducimus. Iure ut sit vitae.", "Nemo optio a unde illo qui. Fugit saepe fugiat molestias rerum qui. Hic et blanditiis aut. Expedita necessitatibus sint ut alias at. Sequi dolores suscipit minus dolor mollitia.", "Asperiores delectus maiores. Porro sapiente accusamus. Rerum voluptas quia earum quaerat autem.", "Cumque necessitatibus laboriosam. Libero perferendis autem itaque. Temporibus autem molestiae omnis adipisci non.", "Eaque ullam deleniti. Omnis aut ut placeat. Consequatur eum est sapiente vitae est ad. Eligendi recusandae excepturi autem culpa. Quae at eligendi consequatur est et ullam ut."]