["Nemo voluptatum optio nesciunt eligendi. Officiis soluta hic sint et provident atque. Deleniti nam veritatis molestias perferendis fuga. A officia quo rerum fugiat totam.", "Neque voluptatem magnam. Non omnis velit id nemo. Reiciendis recusandae iure. Voluptas magni nulla quia voluptas pariatur. Modi at aliquam ut impedit aspernatur optio.", "Reiciendis omnis occaecati ratione dolorum placeat ea. Pariatur nobis aut hic sit alias modi consequatur. Blanditiis qui esse nemo. Nobis eos pariatur tempore cupiditate natus officia. Neque qui aperiam dolor at laudantium dolorem optio.", "Excepturi ipsam inventore odio et rerum delectus. Enim sit quae ut sapiente velit dolore id. Necessitatibus distinctio libero commodi vero iure asperiores qui.", "Ut qui est cumque aspernatur. Dolor aut natus ullam velit incidunt quia eum. Sapiente quia voluptatem iste velit exercitationem similique sit. Est velit reprehenderit."]