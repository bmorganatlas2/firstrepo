["Illo et error mollitia nisi. Aspernatur pariatur vero quis sit qui repellat doloribus. Aut dolorem eaque ea. Eum quas soluta est odio beatae non cum.", "Aliquid quasi consectetur quibusdam. Deleniti temporibus dolore. Quidem consequatur qui.", "Nemo nihil impedit. Qui aliquam quos corrupti aperiam nostrum corporis ipsa. Quae nostrum cum voluptatem ut fugiat ut sed.", "Quis voluptatem molestias illo expedita quod. Alias ipsam neque sit voluptatem similique quaerat. Consequatur autem velit vero voluptatum et cupiditate. Aut minus et.", "Corrupti cumque autem vel nihil. Repudiandae perferendis quia. Maiores soluta commodi sequi et. Sit saepe cum placeat quaerat sed. Sed in accusantium ducimus consectetur tenetur libero."]