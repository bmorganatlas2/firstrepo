["Modi quia beatae voluptatum tenetur. Quia officiis sapiente reprehenderit. Aperiam voluptatem nulla. Voluptatem doloremque exercitationem quas sit.", "At qui nisi aut architecto. Consequatur non quaerat aspernatur ullam tempora eligendi. Et qui voluptas at ut et.", "Natus eum et tempora. Repellendus sint occaecati modi aliquam consequatur. Alias nihil nihil dolore qui.", "Modi dolores sint vero. Qui tempora fugit rem libero nobis officiis commodi. Ut deleniti autem rerum eius temporibus non.", "Aspernatur dolor et. Doloribus in veritatis aliquid error. Vel est consequatur qui eveniet eos dignissimos impedit.", "Laboriosam beatae ut excepturi. Quasi nulla ut debitis unde ipsum omnis necessitatibus. Sunt cumque occaecati optio et laudantium impedit.", "Amet non explicabo voluptas occaecati harum aut. Tenetur ratione sit aspernatur sunt repellat. Qui natus non eos et ut beatae voluptatem.", "Sint doloremque corporis unde vitae consequuntur omnis. Sapiente cumque blanditiis consequuntur dolorum. Incidunt ea vero et.", "Eius inventore velit. Ut cumque tempora. Occaecati quo temporibus et totam non sit. Optio error sed. Iure accusantium vitae."]