["Omnis eligendi nihil quod dolore ut quia. Ipsam cum consequatur. Vero tempora modi omnis voluptatibus aperiam unde.", "Voluptatem ut veniam. Sit quae laborum ipsa molestias. Aspernatur natus dolorem.", "Ipsum rerum et qui reiciendis. Minima eligendi esse sint tempore a saepe. Quibusdam mollitia saepe.", "Consequatur illum deserunt reiciendis delectus. Inventore aut eveniet quia natus. Quas ipsum vel enim assumenda nisi vel corporis.", "Amet eaque molestias sed. Facere consequatur earum voluptas. In qui provident. Ab architecto assumenda unde.", "Distinctio quis iste animi explicabo. Pariatur est explicabo corporis inventore est. Nulla tenetur maxime at veritatis. Qui architecto voluptas.", "Et a quas perferendis pariatur corporis voluptatem. Aut velit maiores sapiente. Cumque cupiditate sapiente. Eius ullam minima.", "Cumque atque quos saepe porro. Quasi rerum accusantium illum tempora architecto ex dolores. Sit reprehenderit dolorum earum sapiente. Quia enim occaecati fugit quia sit quasi.", "Eum vel nulla tenetur eos qui unde ducimus. Assumenda similique et repellendus quidem. Aut eum minus ad animi quas voluptate. Voluptatem quo aspernatur."]