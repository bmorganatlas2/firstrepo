["Voluptatibus similique reprehenderit cumque repellendus. Alias ea fugit. Dolorum est ipsam illo ut omnis. Ut qui sapiente consectetur. Possimus sint quia illo libero.", "Ut saepe dolor. Sit eos ut voluptatibus ut quis saepe. Rerum consectetur sint voluptatem vero. Maiores magni voluptatem.", "Molestiae culpa sint possimus sapiente. Nulla commodi amet nihil nostrum. Quia nihil eum reprehenderit optio atque molestiae. Animi et omnis est voluptates porro dolor.", "Nihil ut magni labore ipsa fuga. Non et veniam. Doloremque accusamus velit iusto nihil id voluptatem tempora. Quidem deleniti placeat. Laudantium voluptatibus quia amet perferendis voluptas at accusantium.", "Cumque et sunt. Saepe minima explicabo. Nemo accusantium omnis ut tempora fuga quis doloribus. Distinctio eaque ratione dignissimos ut sint.", "Quia autem quos qui nemo perferendis et eligendi. Laborum temporibus occaecati omnis. Totam labore veniam qui. Voluptates a sapiente sit ratione quis."]