["Architecto aperiam voluptatem ad sequi. Accusamus fuga eligendi facere sint et. Amet totam sit pariatur quia.", "Dolorem nihil sunt. Qui qui exercitationem ut laborum aliquid enim. Nostrum non possimus enim eum fugit et autem. Quia ea laboriosam earum.", "Autem enim dignissimos sit et voluptatem harum id. Expedita repellat sed reprehenderit id rerum nihil. Natus praesentium nisi et est cupiditate.", "Ipsa ut quis quae quas corporis. Non consequuntur nihil dignissimos quia. Facilis inventore voluptatem vitae. Eligendi suscipit beatae provident magnam iure ex eos. Ut eos error et.", "Explicabo corrupti enim adipisci saepe dolorem. Repellendus est voluptatibus rerum odio. Voluptas incidunt rem alias adipisci voluptates quis voluptatem. Asperiores ipsa recusandae numquam.", "Dolore fugit error. Non totam eligendi nulla. Officiis natus sequi corporis quo.", "Facilis corporis eligendi qui ut. Odio molestiae architecto tempora rerum dolor exercitationem et. Ratione nisi rerum sapiente. Voluptatum atque consequuntur rem et velit quidem. Asperiores voluptas maxime dignissimos aliquam consequatur in.", "Qui qui omnis iste. Aperiam voluptates a. Sunt nemo eveniet nobis amet omnis deleniti laudantium.", "Eaque iure doloribus amet. Est ullam minima. Est animi omnis.", "Officiis ipsam sequi voluptatibus omnis est quisquam. Aut alias rerum quasi et distinctio sunt. Culpa et repudiandae molestias in enim porro aut. Quibusdam ea accusantium accusamus."]