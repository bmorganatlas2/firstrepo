["Et dicta quia. Culpa voluptatem sint adipisci itaque. Corporis et eligendi a.", "Animi ut sunt non soluta. Sint voluptas qui omnis ut. Est qui quisquam. Amet velit dignissimos error explicabo vel est fugit. Vel aut consequatur autem reiciendis deleniti facilis dolores.", "Cum hic quaerat. Sapiente cumque aut occaecati soluta velit exercitationem atque. Adipisci ipsum earum. Provident adipisci quis id animi.", "Culpa officiis quia atque. Tempore nam modi quae corrupti adipisci laborum voluptatem. Laboriosam perferendis quidem reprehenderit aliquid. Error dolorem soluta voluptatem exercitationem. Tempore harum asperiores tempora."]