["Dignissimos dolorem at minima illo et et. Praesentium quidem esse ut quia. Iusto ut et. Deleniti consequatur et quia explicabo ex aut ipsam.", "Rem qui architecto. Cum sit quia soluta. Saepe et earum officia consequatur."]