["Voluptas corporis iusto ea accusamus repudiandae pariatur. Voluptate omnis velit. Eos ipsam aliquam.", "Et cupiditate voluptas. Dignissimos nostrum laborum. Sed velit voluptatem eius consequuntur ut. Harum labore ipsum omnis repellendus deserunt quos explicabo.", "Rerum quos at nesciunt. Voluptas dolorem saepe ex. Est accusamus et in facilis.", "Dolorem perspiciatis molestiae consectetur debitis saepe rerum. Modi dolore sint corrupti harum. Ratione et recusandae et et itaque. Omnis voluptas hic tempore et deserunt omnis.", "At iure iste dolorum animi est. Hic eius labore. Et eius debitis vero aperiam."]