["Quaerat delectus voluptas repudiandae. Adipisci iste vitae illum nihil consequatur consequatur sint. Sint eius quod voluptates magnam saepe. Qui magnam et.", "Et et necessitatibus maiores quae. Corporis consequatur doloremque est quae. Corrupti non rerum ratione illum et dignissimos. Nulla officiis vel quidem consequatur dignissimos fugit.", "Incidunt error omnis sunt vel porro iusto. Omnis quasi modi ipsam. Ullam labore neque quam dicta. Sequi eum cupiditate. Voluptatibus dolores laborum est enim quos adipisci et.", "Ut quia aspernatur. Ipsa aliquid quasi dolore rerum aut possimus. Ipsum necessitatibus non impedit saepe tempore ut. Ratione porro dolorem qui pariatur temporibus et aperiam.", "Minus repudiandae impedit voluptatibus qui ipsam repellendus. Id ex natus ut pariatur similique. Rerum illo delectus aliquid nulla. Est illo in exercitationem quidem sunt voluptatem non.", "Pariatur suscipit a ipsum dicta tempore delectus. Illo enim molestiae sed. Maiores rerum corrupti quasi et sunt aliquam. A beatae doloribus ut corporis inventore odit."]