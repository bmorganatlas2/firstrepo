["Quia error totam nisi est aut aut. Neque ut laborum dolores nihil maxime laudantium sit. Qui voluptas exercitationem ut labore sit.", "Quasi deleniti ut quis. Omnis fugiat corrupti cumque eum delectus impedit. Nisi autem expedita. Voluptatem earum eveniet tempore rerum voluptatem perspiciatis. Quasi non eius.", "Animi maxime optio voluptas tempore unde veritatis asperiores. Error dignissimos incidunt quo exercitationem reiciendis. Voluptatem quaerat dolor et consectetur et.", "Laboriosam rerum dolor eius quia. Illo fuga tempora voluptatibus ut. Reiciendis deleniti tempora porro minima at quia excepturi. Molestiae laudantium pariatur corrupti. Aut dolorem sunt qui totam qui."]