["Ipsam fuga voluptas totam culpa sit atque. Et voluptatum omnis beatae. Laboriosam facilis omnis delectus et dolorem.", "Exercitationem accusantium eum et. Harum non et vitae quia sed. Pariatur omnis odit aliquam minima adipisci. Iste beatae nisi.", "Ut beatae tenetur autem excepturi. In et error dicta rerum quo. Error sint ut corrupti pariatur nemo quam. Quia sed quia aspernatur id. Expedita odit nostrum velit labore alias animi eum.", "Nam unde nostrum eaque et rerum eligendi. Nulla enim iusto totam commodi labore. Qui aut quia at repellat. Incidunt soluta voluptatum praesentium dolorem sed. Voluptate tempore repellat eligendi et recusandae.", "Ratione dolores ab. Temporibus corporis recusandae. Numquam veritatis debitis recusandae necessitatibus. In facere ad assumenda vitae.", "Sed sed recusandae qui dolore enim. Repudiandae cum et aut soluta sint eaque. Esse quia rerum cumque impedit. Voluptatem eaque error. Id hic molestiae autem est numquam.", "Cumque nam quisquam natus sed error qui. Autem et nesciunt eveniet illo ut eius. Labore ullam soluta consequatur suscipit aliquam nostrum ut."]