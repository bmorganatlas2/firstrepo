["Quia quo incidunt vitae laborum rem et corrupti. In eligendi ipsam ut omnis iste ab ut. Veniam aut porro velit ea quia ut qui. Error ipsa molestias sit voluptas.", "Eligendi consequatur velit optio facilis qui vel impedit. Optio sint debitis aliquid asperiores molestias nobis amet. Veritatis delectus dolor non.", "Aut esse dolores ducimus ipsum magnam modi et. Velit hic voluptas voluptatem. Voluptates minus neque quia mollitia consequatur facilis.", "Necessitatibus qui eligendi corporis explicabo. Dolore rerum at vitae doloribus voluptatem sunt. Qui maxime a dolor fuga. Eos exercitationem dicta dolores.", "Sed odio est consequatur est harum voluptatem. Sed laudantium vitae eveniet. Est et voluptatem atque consequatur sed quaerat voluptas. Voluptatibus et reprehenderit est et.", "Sint incidunt corrupti nemo officia quia. Amet iste quo esse tempora. Aut quia mollitia nostrum dicta quo."]