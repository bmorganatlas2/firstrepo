["Ipsa quo qui earum sunt. Dolores excepturi exercitationem ad labore ut placeat et. Aspernatur aliquam id quisquam sed autem repellat quia. Rem doloribus facere iste dolores molestiae laudantium sapiente."]