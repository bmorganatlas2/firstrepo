["Qui id officiis. Aut ipsum aut temporibus eaque ea itaque. Sunt numquam ut repudiandae illum.", "Sed eum inventore repellat et omnis. Aspernatur eos illo et. Similique fugit doloribus voluptatibus.", "Quod fuga assumenda quis cum. Nobis dolores iste. Aut repellendus dolorem necessitatibus. Corporis error odio omnis eos reiciendis ut repellendus.", "Necessitatibus et qui amet est enim dolor officiis. Dolores ut eaque aut laudantium laboriosam. Nemo beatae at optio aliquam molestiae. Quia maiores omnis ab eum dicta nostrum dignissimos.", "Eum sit recusandae. Neque dolores odit aspernatur qui. Velit voluptatum minima et doloremque consequatur veritatis. Aliquid qui cupiditate doloremque nostrum assumenda est. Quia voluptatem eveniet omnis.", "Ratione alias rerum minima et. Est repellendus quia architecto quos magnam maiores dolorem. Ipsa quas et exercitationem dolorum nostrum quos laboriosam. Laudantium cumque iure.", "Maiores aut qui. Rem quo doloremque soluta vel ut iste dolorem. Nesciunt quos repudiandae. Accusamus voluptatem nihil nam sint sit non velit.", "Quidem omnis voluptate atque. Quam inventore qui molestiae. Perferendis laborum sint consequatur eos debitis non autem. Velit corrupti adipisci. Nulla quia voluptatem natus doloremque tempore eaque possimus."]