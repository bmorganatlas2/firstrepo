["Earum deserunt neque necessitatibus optio veniam quo ipsa. Perferendis ex et aliquam. Perspiciatis placeat similique aut eos quis. Necessitatibus odio expedita neque et provident ea doloremque.", "Laboriosam rerum voluptatem ullam optio laudantium dolores et. Ipsam quia aperiam qui ex ratione. Et perspiciatis ex. Voluptatibus unde amet.", "Consectetur rerum cum qui iste dolores quod. Nulla voluptatem dolorum optio quisquam cumque. Dolorem praesentium voluptatum voluptas qui.", "Harum eveniet veniam id magni aliquid atque. Esse itaque et. Et in non. Rerum eum architecto mollitia sed explicabo.", "Nulla iste error doloremque in eveniet qui fuga. Ut similique veniam quidem laboriosam earum. Sit eos laborum.", "Est architecto labore blanditiis iusto. Repudiandae omnis sed enim. Iure natus sunt unde tempore. Aut qui quis mollitia quia qui non animi.", "Illum iusto inventore aliquid sint exercitationem. Et exercitationem voluptatum incidunt quo maxime non perferendis. Aut quibusdam quis. Mollitia eos est delectus dicta sequi odit perferendis. Nihil voluptatibus veniam temporibus nulla libero.", "Et et ex odio deleniti. Qui sit magnam. Laudantium nam ipsam. Et sint et quae."]