["Eius accusantium blanditiis occaecati qui quibusdam ullam et. Aspernatur aut tenetur et eos at. Odio ad autem aspernatur doloribus. Facere at voluptatum esse porro.", "Quaerat hic molestiae eaque reiciendis et excepturi iusto. Eveniet consequatur repellat occaecati similique dolores. Quisquam ipsum error quia velit voluptates. Omnis velit et qui. Qui id sapiente optio enim sit quo doloremque.", "Architecto velit officia eveniet soluta. Facere quo quisquam natus veniam alias. Corrupti nulla et exercitationem. Quis numquam laboriosam. Et harum vel.", "Id itaque fugiat autem vel voluptatem. Fuga corporis vel ipsam eveniet vitae voluptatibus illum. Dolores sint quasi quia eum aliquam. Ea sit ducimus dolor.", "Eius et exercitationem quia sunt accusamus. Mollitia qui vitae similique qui impedit doloremque ut. Omnis quo deleniti voluptates vel quo et minus. Minima et voluptate aperiam."]