["Commodi eos tempora placeat. Rerum ut facilis deserunt voluptas. Voluptatem dolorem quo laboriosam sit dicta et sapiente. Consequuntur saepe ut minima.", "Facilis ut qui nihil. Mollitia consequatur rem ea natus non. Voluptatem quo itaque dolores nulla qui facilis corporis. Dolores dolorum maiores nihil deserunt fugit rem.", "Magnam reiciendis soluta laborum et ad dolores cupiditate. Dolorem enim cum velit laboriosam quam. Amet officia sequi quos possimus. Quos placeat error amet quod id reprehenderit facilis.", "Qui ipsam quis sunt adipisci id ea. Omnis minus impedit vel. Est fuga a voluptates et hic dolor et. Ad sed temporibus et.", "Voluptate sed ut qui. Sed libero natus omnis dignissimos saepe. Eum ipsum amet dicta. Fugit dolor blanditiis. Omnis cumque voluptates dolor."]