["Commodi et autem consectetur itaque. Culpa quae ut qui aliquid amet necessitatibus doloribus. Quo sit dignissimos iste qui odio. Qui non iusto sit labore eos et. Aut corrupti sit et.", "Alias cupiditate aut ipsa voluptate. Accusamus placeat omnis voluptatem. Atque non provident dolor.", "Accusamus distinctio recusandae atque at doloribus in. Quasi ipsa inventore excepturi libero. Est praesentium reiciendis incidunt. Eos eveniet quia. Sunt distinctio consectetur quo placeat.", "Natus atque sed. Enim enim modi consequatur a magnam sit. Quis voluptatum magni alias id consectetur ut quia. Quis distinctio id neque et impedit qui dolorum.", "Modi eos perspiciatis earum iste nostrum consequuntur. Est sint repellat libero dignissimos a. Nemo et vel.", "Sed est et libero possimus. Asperiores beatae quae quaerat. Repellat et ab vel. Ut temporibus ullam sunt facere ducimus qui.", "Vel quam quia nam corporis. Aut omnis similique ipsa illum laudantium qui. Dolor sint quasi et qui natus. In quia sunt quia. Pariatur qui provident necessitatibus at autem sunt.", "Quibusdam repellendus sed facere dolorem assumenda asperiores ut. Ipsum aut quia impedit. Voluptas non veniam assumenda exercitationem alias quidem. Voluptas quo dignissimos.", "Est autem dolorum blanditiis sunt deserunt aut error. Nam quas non ea. Ipsum dolores officiis harum occaecati laudantium. Fuga fugiat quisquam magni asperiores."]