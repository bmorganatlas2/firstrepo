["Qui expedita rem sed pariatur vel minus. Dolores assumenda voluptas odio aut fuga laboriosam expedita. Accusamus in nostrum qui porro ea. Eius est quis neque earum animi dolorum occaecati.", "Animi sed omnis accusamus est. Adipisci incidunt qui facere esse fugiat molestiae optio. Rerum blanditiis est porro vel est sint laudantium. Aliquid impedit voluptatibus quo quia rerum.", "Cumque quas eveniet. Hic est rerum aliquam alias quaerat omnis eveniet. Rerum quaerat dolores veniam iste ducimus ut. Illo illum voluptatem a sint minus.", "Qui non neque. Molestiae impedit eius quis accusantium temporibus vel. Possimus sapiente quisquam fugit delectus consequatur perspiciatis.", "Deserunt odit quisquam sapiente enim pariatur. Consequatur voluptatum ipsam sequi. Rerum qui quia dolorum explicabo ea adipisci. Quo sed incidunt voluptatum quis. Autem nostrum voluptas.", "Eum odio aut consectetur. Aliquam suscipit asperiores nesciunt nobis quod ut deleniti. Qui consequatur aut minima nemo quaerat.", "Qui quasi praesentium quidem accusantium. Cupiditate id nemo praesentium non reprehenderit. Alias reiciendis doloribus ipsa unde qui. Enim molestiae earum. Sint incidunt molestiae cupiditate.", "Et occaecati amet ex quae qui voluptates cupiditate. Non perspiciatis cupiditate. Atque ullam voluptatem.", "Voluptatum quo sit explicabo. Neque est harum atque sit delectus autem. Est impedit temporibus sit nisi architecto. Unde impedit vel assumenda. Aut est temporibus porro sed dignissimos in.", "Possimus accusamus sit et earum culpa. Harum eligendi doloremque libero ut perspiciatis corporis asperiores. Qui qui omnis ipsa est. Voluptatibus veritatis dolores possimus excepturi."]