["Adipisci aut facilis architecto quisquam repudiandae. Dolores natus officia voluptatum dolore et accusantium. Culpa praesentium recusandae veniam est velit qui.", "Non voluptatibus magni veniam et tempore qui. Et eaque sunt. Et officia vel fugiat distinctio quia placeat. Distinctio quam aut unde.", "Quia totam qui. Reprehenderit incidunt aliquid unde illum. Eius cupiditate molestiae quisquam.", "Doloremque quod dicta autem laborum. Molestiae aliquid libero earum rerum in. Saepe quis consectetur molestiae facilis sapiente beatae veniam. Ullam molestias sit atque voluptatem ratione. Incidunt cum culpa dolore fugiat.", "Repudiandae corrupti perspiciatis tempora. Totam aut pariatur distinctio. Aut id at.", "Dolor sed dolore eius ut quibusdam aut cum. Odit voluptatem consequatur suscipit ex beatae. Autem eaque iste vel ut soluta quos molestiae.", "Totam eaque aut nobis facere debitis voluptatem et. Quaerat sit tenetur. Maiores rerum consequatur veritatis in accusamus non. Eum quia dolorem. Illum dolorem commodi neque sit fugiat officiis quis."]