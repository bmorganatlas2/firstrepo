["Aut voluptas quo asperiores alias. Similique reiciendis consectetur officia. Saepe ut accusamus nihil suscipit tempora fugiat a. Praesentium esse quae a officia rerum earum hic. Maiores nisi magnam.", "Ut est dolorem omnis quos id hic. Velit qui eos est possimus id consequatur autem. Incidunt laudantium blanditiis distinctio sit. Aut excepturi qui aperiam amet laborum officia incidunt.", "Voluptatum voluptatibus nam aperiam odit. Pariatur sint hic et quidem dolor nesciunt voluptates. Sed quis voluptas atque. Quae beatae doloribus neque fugiat ad voluptatem labore.", "Soluta quod unde voluptas. Tempora itaque et totam beatae excepturi. Est non molestiae cupiditate quia et similique rerum. Voluptatem ut labore similique iste temporibus facere. Quasi ea ut aut in officia.", "Ut quia ut et reiciendis. Consequatur tempora nesciunt optio laudantium accusamus fuga eos. Odio consequatur esse culpa facere tenetur.", "Ex omnis eveniet dolore ipsa. Culpa voluptatem magni blanditiis occaecati est. Et debitis corrupti saepe labore mollitia quos voluptas.", "Suscipit odio ut. Laborum ab eum quia rerum et cum. Dignissimos distinctio dolores rerum similique doloremque beatae sint. Fugit ea cum debitis accusamus. Et velit dolor.", "Ut nihil aut omnis. Nam vero non. Iure impedit velit repellendus nostrum explicabo ducimus maxime.", "Vitae nam atque corporis. Officia ut aliquid aut labore dignissimos. Autem excepturi rerum officiis quae ullam sunt. Animi voluptas sunt reprehenderit in harum commodi nihil."]