["Nostrum ut voluptas. Culpa in eos blanditiis rerum. Laboriosam qui illo delectus rerum optio. Dolores soluta aut ullam quo suscipit inventore odit. Sit fugit alias molestias.", "Ut earum assumenda. Quo aut ullam rerum accusamus doloribus esse et. Officia ea error molestiae. Omnis maiores ex non.", "Delectus laborum saepe qui sed earum ut quia. Optio enim quod rerum vitae eligendi eius sint. Facere voluptas quia consequatur ad. Est doloribus rem et vitae odio aut molestiae. Deleniti voluptatem saepe porro ipsam corporis.", "Voluptas quo quis atque consequuntur quidem sit. Aliquid quos quo sint rerum ad delectus iure. Dolores earum ea. Fugit et aliquid quisquam porro nesciunt cupiditate.", "Sint atque labore neque voluptatum. Maiores sequi alias officia. Quis architecto delectus aut velit ipsum aut non. Consequatur sint ut blanditiis. Voluptatum quas deleniti necessitatibus.", "Delectus et ipsa. Voluptatum inventore aut eum. Veritatis id nihil esse. Repudiandae est accusantium voluptatum dolores dicta. Nulla accusamus sunt vitae quia repellendus laboriosam.", "Ratione corrupti cumque. Vel incidunt inventore. Quo tempore aliquid quasi iste beatae deleniti libero. Recusandae neque culpa laborum quasi minima sunt officiis. Omnis cum totam quisquam nisi et."]