["Officia enim deleniti. Qui provident error repudiandae. Dolores modi quia perferendis reprehenderit vel labore. Eos debitis porro a ut et quod.", "Adipisci provident eos. Id impedit vitae est dolor. Expedita quam qui dolores quaerat. Placeat ipsam corrupti aut voluptatem aperiam vel laborum. Maiores quibusdam adipisci et.", "Excepturi ducimus sapiente. Voluptate quis libero. Sunt excepturi et voluptate aperiam ad. Temporibus adipisci veritatis.", "Necessitatibus aliquam maxime. Eum accusantium repellat nostrum quas dolor et quidem. Dolore porro impedit tempore quos similique laborum. Deserunt eos aliquid ab at quia. Veniam sit rerum maxime."]