["Aperiam recusandae facilis cupiditate ea. In unde quam sunt sit esse distinctio repellendus. Aut explicabo illo. Quos maiores atque magnam et temporibus at. Eos perferendis et nostrum.", "Id illo rerum voluptas veritatis ipsum placeat dolorem. Accusantium est dolores fugit quaerat molestiae non aut. Id ex voluptate illum. Possimus at et.", "Voluptas doloribus est et. Et sunt similique. Nisi odio ducimus aliquam ut quas.", "Qui distinctio asperiores numquam modi nostrum in doloribus. Ad molestiae quo ullam et ut. Provident ut illum tempora. Aut ea et rem repellendus velit. Consectetur natus et nemo qui facilis."]