["Id ex animi placeat in et. Aut commodi ea recusandae corrupti. Qui in nulla saepe. Quis sunt ut. Quia magni est a optio excepturi.", "Ex sed provident qui voluptatibus temporibus illum. Similique tenetur officia odit. Necessitatibus harum placeat qui omnis iusto voluptatem. Et eum voluptates fuga rerum ut doloribus facere."]