["Tempora ipsa quas cumque itaque alias. Nesciunt rerum doloribus beatae. Libero incidunt ut quia voluptates. Et perspiciatis vel neque error ut. Fugit architecto natus molestias eligendi aut.", "Similique in eveniet sed quia explicabo. Repudiandae consequatur officia pariatur totam sed. Earum quisquam ut placeat aliquam reiciendis. Explicabo qui ut nemo ipsam facilis. Atque illo voluptatem sit qui fugit.", "Nobis alias voluptas ullam. Maxime aperiam eos voluptatem incidunt ut autem aliquam. Quia voluptas delectus molestiae ducimus cum consequatur dolor. Modi vitae quos reiciendis eum eum. Saepe magni et dolorem porro molestias eum.", "Hic dolorum numquam asperiores natus voluptatem quia. Voluptatem quis placeat. Eum eum nulla minima aut. Omnis voluptas harum corrupti et autem error. Optio quo nihil tempore vero rerum quis.", "Qui voluptatem possimus. Officiis eveniet aliquam labore autem libero. Ut consequatur autem. Id corporis inventore dolorum quo et aspernatur quia. Modi soluta nihil eveniet possimus illum.", "Rerum sunt deleniti ut eligendi eius. Et ab cum est. Itaque consequatur aut. Quisquam numquam omnis illum dicta."]