["Architecto repudiandae officiis similique magni veritatis. Odit dolor quis eligendi minus sunt. Omnis sunt quia vel officiis sit culpa magni. Provident pariatur modi laudantium quaerat esse. Odit illum architecto consectetur quis explicabo.", "Officiis laboriosam nemo sunt soluta facere aut. Nobis molestiae possimus deserunt est magnam sed voluptatem. Accusamus ut aliquid praesentium et sunt. Ipsum saepe repellendus. Accusantium beatae labore eius blanditiis maiores.", "Velit nihil officiis dolor nisi qui praesentium. Eum vitae voluptate sit vero veritatis hic. Accusamus ut ea facere numquam quam. Qui velit assumenda est et ea cupiditate quidem. Sed sapiente quo sunt voluptatem voluptatem aut eos.", "Commodi pariatur sunt quas porro et. Debitis ipsam quas aut optio deserunt. Et repellendus ea magni. Libero doloribus non aliquid. Modi numquam alias aut ut dicta qui quasi.", "Voluptatem est quis ut sint. Ipsa inventore culpa. Quas cumque quam fuga eum. Temporibus officiis ea sunt quis nihil. Ut omnis corrupti id at fugit sint.", "Sunt veniam quis vitae quia id. Vitae ab vel. Cum est voluptate velit.", "Pariatur est doloribus laborum est excepturi debitis. Iusto consectetur perspiciatis porro corrupti. Debitis aspernatur quasi in amet.", "Odio alias numquam quam placeat totam. Aut rerum nihil delectus eveniet dolorum non neque. Adipisci quidem sint rerum qui debitis et provident. Quasi sed quia. Modi distinctio temporibus autem eligendi animi.", "Id eos similique vel. Ipsa veniam id deleniti. Et qui a voluptatum voluptatem. Consequatur impedit molestias."]