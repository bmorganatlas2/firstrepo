["Quae molestiae commodi. Autem exercitationem qui adipisci omnis iusto quos voluptatum. Quo sit repellat consequatur vero voluptate.", "Totam quam commodi cumque quia animi. Repellendus quo provident. Sunt dolor aut quia enim harum illo reiciendis. Non sed nulla accusantium qui minus.", "Quod aperiam repudiandae laborum dolore provident quo. Dolore rerum vitae recusandae. Minima commodi facilis voluptas.", "Modi unde doloremque laborum magni aperiam fuga odio. Est aut enim consequuntur minima laudantium. Ad deleniti magnam eius nam quae maxime ratione.", "Cupiditate quia rerum corrupti hic ducimus. Dignissimos recusandae ut. Provident ea rerum voluptatem quod molestiae est. Rerum et consequatur amet minus.", "Ipsa odio exercitationem. Necessitatibus deserunt eius. Consequatur consectetur provident."]