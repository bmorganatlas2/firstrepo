["Est ut reprehenderit consequatur quia aliquam voluptates laudantium. Quo quia dignissimos possimus placeat dolor. Eligendi laudantium officiis dolores. Necessitatibus omnis natus.", "Voluptate quaerat enim dolor id. Beatae architecto possimus enim cum autem aut voluptas. Dolore iure voluptate quia.", "Nostrum atque voluptate temporibus dignissimos nemo quae. Voluptates nihil voluptas provident. Beatae ducimus voluptatem.", "Vel rerum molestias mollitia perferendis similique officia. Molestiae earum tenetur aut sunt. Natus dolorem dignissimos repellat ratione est quasi reprehenderit. Nulla alias et maxime et ut.", "Ex eius vel. Quasi fuga et qui possimus enim in. Iusto neque sit est adipisci et. Libero nihil repellendus assumenda maiores."]