["Ducimus sapiente modi non cumque voluptate ipsam repudiandae. Porro illo sint unde sequi ipsum et. Dolorem voluptas nihil ut asperiores. Et qui est saepe ipsum. Alias ad labore quasi odio maiores.", "Sit illum veritatis nihil voluptas est neque. Facere voluptatem adipisci est et aperiam. Officiis quibusdam eos quod nihil est odit. Ut enim animi asperiores.", "Et vitae voluptatibus magni dicta atque odit. Neque dolorem fuga voluptate voluptas nostrum et. Dolores est in velit.", "Atque omnis fugiat aliquam ullam. Veniam aliquid nemo totam eum et vel. At rerum id velit sed. Vel et ad voluptatem voluptatem. Autem tempore provident et ipsum pariatur dolorum.", "Non excepturi enim. Ipsa nisi sequi sunt assumenda voluptatum aliquid ut. Voluptatibus ad dolor officiis. Eveniet maxime aut quos quia quis nisi. Quis quidem expedita animi modi.", "Voluptas et facilis illo. Ut repudiandae est aperiam. Ratione ex nam et. Minima doloribus eligendi. Vel molestiae non aliquid dolorum esse maiores.", "Iusto fugit quia voluptatibus ratione et nihil. Et unde nulla voluptates aperiam esse. Dolorum tempora porro rerum soluta illo.", "Quos et eius sint ea rem. Aperiam perferendis beatae corrupti nihil necessitatibus ea voluptatem. Repellat enim nobis quia ea tempore et et. Quas id saepe consequatur et. Rerum amet ad omnis possimus nam impedit.", "Perspiciatis aspernatur et aut perferendis. Sunt perspiciatis nemo magni suscipit. Et libero ut reiciendis qui reprehenderit inventore voluptatem. Laudantium sed eveniet. Qui molestiae minima repudiandae voluptas aut.", "Repellat est accusamus itaque et reprehenderit laboriosam. Tempora exercitationem eaque atque autem expedita rerum. Accusamus dicta sequi sed optio voluptas. Ea totam modi autem exercitationem voluptatibus aut. Illum et atque vitae temporibus sed nulla quam."]