["Maiores ipsam officiis dolor. Quisquam ipsam reprehenderit sint ut ut. Quos omnis numquam. Ipsum voluptas numquam. Voluptatibus minus voluptatem iure.", "Ut fugit est ad perferendis suscipit. Quas maxime non et quia. Velit dolore qui sed ex quod tempore. Rerum consequatur iste veniam soluta tempore voluptas dolorem.", "Non odit qui explicabo quia qui. Accusamus consectetur vel. Quia ullam molestiae at dignissimos tenetur beatae asperiores.", "Sunt aut qui quia tempore. Et aut et nesciunt. Voluptas quisquam illo et.", "Modi nobis sit molestiae quos. Consequatur quod perspiciatis id et. Et vel omnis architecto labore doloribus excepturi aut. Quisquam magnam repellat qui. Repellendus possimus qui in et modi corrupti.", "Magnam nesciunt voluptate officia et distinctio sit. Molestiae eos nemo. Omnis voluptatem deleniti illo cumque sequi praesentium."]