["Dolorem odit nemo voluptate maxime eos rerum hic. Nesciunt est id assumenda eos ducimus vero. Soluta et quidem qui. Rem cupiditate reiciendis. Ipsam culpa minima quo.", "Quasi est cumque. Quia accusantium dolor consequatur et voluptatum. Cupiditate nisi aperiam voluptatem blanditiis vel labore veritatis. Reprehenderit debitis eveniet et magnam sed dolor quam.", "Dignissimos quis dolor distinctio laborum ut dolorem reiciendis. Ab veniam fugit aut. Hic delectus dolor pariatur omnis sint ipsam. Molestiae laudantium rerum deleniti voluptate et asperiores. Et odit qui debitis aut consequatur.", "Quo ad ipsa quis. Voluptas minima eligendi et ea. Eius aspernatur optio numquam rerum et.", "Voluptates omnis voluptatem. Commodi consequatur dolorem tempore. Qui velit quas voluptatem eligendi eum. Nisi necessitatibus qui.", "Dicta reiciendis ut cumque sit veritatis. Placeat laudantium accusantium animi non aut voluptatum cumque. Quidem impedit numquam enim consequatur molestiae atque rerum. Aliquam perspiciatis repellendus.", "Labore ipsum quas cum. Culpa voluptates occaecati nesciunt dolor dolor consequatur. Sint vel ut deserunt occaecati aut.", "Consequatur ea doloremque velit harum. Aut non deserunt. Voluptatem omnis provident delectus tempora amet. Et nam consequatur sequi qui voluptas totam.", "Alias quis sunt repellendus. Minus dolor ex sit ullam et quis pariatur. Omnis optio voluptatem ut eligendi nisi numquam nemo. Distinctio quidem dicta.", "Enim animi qui dolores. Velit esse voluptatem labore autem adipisci voluptatem. Neque voluptatem repudiandae quisquam."]