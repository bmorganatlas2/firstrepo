["Corrupti ea qui rerum dolorum itaque voluptas. Dolores reprehenderit in. Iste velit ut tempore doloremque. Voluptatem assumenda molestiae ab harum expedita exercitationem illo.", "Sunt eius porro expedita facilis vel. Dolore doloremque provident. Sint illo adipisci fugiat est dicta vel. Ipsum eum aut. Tenetur sapiente reiciendis necessitatibus dolore qui amet.", "Quisquam harum dicta quibusdam perspiciatis adipisci. Ut consequuntur consequatur eum provident sed qui. Libero et unde rem molestiae. Porro voluptatem dolores saepe cum.", "Sapiente qui veniam voluptatibus perferendis qui. A quaerat consequuntur velit. Nesciunt ut voluptatem. Ratione voluptas adipisci rerum.", "Rerum sequi assumenda est ad ullam laborum. Ipsa necessitatibus aspernatur et molestiae eos. Veniam et eum repellat. Sapiente et omnis aut suscipit. Necessitatibus omnis ut nesciunt eius reprehenderit facilis.", "Est voluptate voluptatem. Est pariatur dolores. Aut quaerat magnam explicabo atque similique consequatur. Eius dolores inventore nesciunt qui eos rerum in."]