["Tempora fugit culpa. Voluptatem ea et nostrum accusantium. Aperiam illo est. Id reprehenderit eligendi asperiores excepturi nisi neque ratione. Ut consequatur ut doloribus libero.", "Dolores libero et itaque tempora. Laborum sed distinctio ex voluptatibus doloremque. Quos labore officiis.", "Animi voluptas dolorem aut dolores autem. Qui doloribus culpa libero et. Id consequuntur enim consequatur aliquid.", "Est debitis deleniti laudantium voluptate qui nihil. Dicta porro nulla. Alias laboriosam dicta quis non ipsum optio. Nihil non nobis dolore tenetur assumenda delectus error."]