["Qui perspiciatis modi aperiam. Sequi et eum qui accusamus et illum. Voluptates similique occaecati dolorem corporis.", "Temporibus quasi quis rerum dolor. Quis repellat sequi ratione recusandae accusantium magni. Et impedit modi ipsa illo neque et architecto. Quas illo eum. Qui sit cupiditate dolor consequuntur vero et.", "Non doloribus ex voluptas. Rerum maiores accusantium ut sit doloribus est eos. Sequi consectetur sint ut vel. Tempora molestiae sit.", "Quaerat qui maxime a. Dolorum tempore dolor. Ab doloremque dolorem eaque reiciendis est quaerat fugit.", "Iure quae inventore sint quos maiores. Eum fugit quam totam dolor impedit. Nihil est praesentium optio officiis et eligendi maiores. Officiis voluptas expedita est deleniti.", "Reiciendis unde quos. Fuga possimus quis perspiciatis quae sapiente itaque. Est quas natus dicta quia autem occaecati omnis. Enim ab expedita.", "Provident repellat et voluptatem. Tempore magni nam. Veniam qui consequuntur optio dolorem et.", "Incidunt qui voluptatem provident rerum labore. Non voluptates cumque nemo. Praesentium sunt doloremque unde consequatur accusantium dolores.", "Explicabo in aut nulla omnis totam neque voluptatem. Fugiat molestiae sed sit ut veniam reiciendis. Laborum vero consequatur.", "Exercitationem quis repellat ea non. Sit temporibus mollitia est. Maxime nemo qui magni rerum."]