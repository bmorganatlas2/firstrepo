["Non est earum ut nulla quas deserunt similique. Laboriosam laborum autem nam. Est et rerum quam non similique exercitationem. Reiciendis illo suscipit impedit. Sint molestiae sapiente ut at.", "Consectetur atque dolorum. Non optio ipsa. Ipsa dolorem quam perspiciatis dolorem laboriosam sed. Aut velit repellat atque voluptas tempore sit. Distinctio harum exercitationem id."]