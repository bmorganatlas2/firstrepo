["Aut repudiandae molestiae quas reprehenderit cupiditate. Omnis fuga et dolor ipsa minima. Accusamus molestias facilis a eveniet temporibus.", "Dolorum delectus rerum aut velit maxime molestias recusandae. Omnis porro ut recusandae consectetur mollitia ab. Minus dolor eius."]