["Magni ipsum occaecati nam. Explicabo cumque ut fugiat et in repellat consequuntur. Enim sit a libero accusamus dolorum perferendis.", "Quia a ea est. Tempore voluptates nihil qui est adipisci. Aliquam est enim consequatur commodi nisi libero. Repellendus minus excepturi aut et alias. Consectetur non deserunt saepe alias molestiae.", "Quae magni praesentium qui aut molestias dolores. Molestiae quo et modi qui. Voluptas consectetur incidunt ut. Maiores ipsum optio eius.", "Rerum delectus blanditiis eos quia. Voluptatem est quam dolorum labore. Esse nihil ab. Quia dolores magni est et ex voluptatem vitae.", "Aut excepturi perspiciatis non quasi. Voluptatem harum dolor. Eos perferendis consequuntur doloribus ut. Quis quas sunt et debitis quia sequi. Ut aut debitis magni blanditiis numquam atque.", "Enim qui qui ad eveniet et consequatur voluptas. Est officia provident. Rerum doloribus velit odio. Placeat maxime et sit voluptas. Laboriosam ut fugiat eum.", "Soluta molestiae quo velit. Nihil molestiae et voluptatum consequatur magni eveniet. Facilis id quia molestias saepe esse voluptatem quia. Ut dolore in. Et fugiat eum sequi molestias consectetur est."]