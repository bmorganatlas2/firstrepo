["Perspiciatis sit officiis omnis asperiores consequatur qui consectetur. Voluptatem accusamus sunt blanditiis. Explicabo sunt tempore eum quos quasi. Dolores voluptatem provident facilis omnis. Consequatur delectus quam.", "Deleniti quo et quisquam. Aut ut necessitatibus ad est rem. Esse voluptatem et quasi. Nostrum iusto autem ea dicta rerum quos quibusdam."]