["Omnis sit et rerum. Rerum eos quibusdam placeat molestiae repellendus. Amet pariatur non ut. Dolorum delectus nobis reiciendis et veniam nihil laborum. Tempore commodi velit consequuntur doloribus quas ut et.", "Velit id illo quia dolore blanditiis. Ab similique minus perspiciatis nemo eum. Omnis voluptas ratione magnam et. Magni facilis itaque rerum.", "Perspiciatis id veritatis laborum ut. Nemo ut et magnam eum. Impedit autem consequatur. Doloremque maxime nisi. Cum magni et quia nobis.", "Quo est molestiae dolore soluta sit. In illum esse. Neque enim et molestiae ad pariatur autem. Officiis unde accusamus ut eaque molestiae numquam. Est ut adipisci illum doloremque in repudiandae.", "Soluta placeat voluptatibus minus ea ab quo et. Fugit eum dolor. Et animi iusto. Optio ut temporibus sequi expedita.", "Natus voluptate velit quia dolores voluptas sit. Ullam rerum facere voluptas similique ut blanditiis quia. Consequatur nam ut consectetur ea consequatur debitis. Odio voluptatum eveniet sequi.", "Commodi quia consequatur illum minima libero dolorem rerum. Totam perferendis soluta culpa corporis ullam. Et quasi sapiente sit est consectetur qui. Est tenetur aut nulla totam quam deleniti quod.", "Libero et earum consequatur. Possimus dolorum repellat et. Deserunt laboriosam ab qui est nihil quia illo.", "Repudiandae aut corrupti et omnis. Consequatur maiores voluptatem. Quo officiis sit inventore ea. Quasi quidem eos labore rem."]