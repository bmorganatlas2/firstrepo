["Autem aspernatur dolorem a nam temporibus qui veritatis. Occaecati cumque et alias in maxime. Quia perferendis ea nobis laudantium consectetur nostrum. Ea vero nesciunt in et quas.", "Occaecati voluptates necessitatibus eos eos voluptatem aspernatur qui. Rerum provident odit facere. Vitae quo perspiciatis nulla.", "Aut alias et ea. Libero illo nihil error vero. Rerum aut quia. Blanditiis incidunt distinctio minus deserunt. Quo repellendus esse eos molestiae.", "Accusantium ipsam fugiat voluptatem dolorum delectus nobis. Doloremque repellat nulla ad reiciendis. Distinctio aut fugiat provident nesciunt modi. Enim vitae iusto quia. Maxime veritatis eum enim consectetur.", "Qui omnis ipsum odio. Fugit accusamus est. Eligendi dolorum iusto laudantium ea voluptatem."]