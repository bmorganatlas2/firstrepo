["Autem qui eius possimus saepe nulla eveniet. Laudantium consectetur non minima odit quae ex. Fugiat et in ullam pariatur et quia dolores. Laudantium quae eligendi temporibus. Voluptatem corporis dolor.", "Incidunt repellendus et quia voluptate earum doloremque deleniti. Et qui in quam. Quam sunt impedit veniam est provident. Culpa non sunt.", "Ducimus sunt expedita iusto nostrum. Laudantium sit quisquam. Odit magnam laboriosam et dicta voluptas aut. Excepturi iste similique possimus debitis quia aut tempore."]