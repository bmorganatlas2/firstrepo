["Nihil ab est omnis aut quia. Qui dignissimos est cumque ratione quia minima. Dolores aut ipsam porro mollitia atque assumenda occaecati.", "Ratione voluptatem qui. Veniam quibusdam labore totam. Officia consequatur sapiente enim rerum reiciendis tempora amet. Autem cupiditate vel.", "Cupiditate magnam eligendi similique. Sequi sit amet et non assumenda qui error. Qui quaerat cupiditate. Perferendis vel est sed magni doloribus. Dolorem tempore dolores illum non unde voluptatem blanditiis.", "Inventore dolor unde. Quia veritatis consequatur aut consectetur ea maxime illo. Et cupiditate nobis et.", "Quia quis similique id velit. Doloribus laudantium rerum occaecati iure accusamus dolorem. Unde dolores voluptatem doloremque nisi omnis voluptas magni. Libero aut non. Eaque itaque quis commodi odit quia.", "Rerum suscipit occaecati quos voluptas autem. Tempora recusandae qui sint laudantium. Aut provident molestias laboriosam quia quia blanditiis occaecati.", "Incidunt distinctio ut praesentium. Explicabo dolorum voluptas eum in voluptatem necessitatibus. Distinctio aut deserunt quia non aspernatur officia est.", "Magnam est perspiciatis rerum id quam. Cumque autem nihil minus debitis. Sit modi doloribus molestiae omnis est fugiat minus.", "Nam laudantium tempora est cupiditate molestias. Consequatur voluptate molestiae magnam voluptatum similique est in. Voluptas ut totam neque praesentium rerum facere. Ab et ea."]