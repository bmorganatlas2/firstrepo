["Ad quo qui autem tempore porro et ab. Hic cumque minus. Non temporibus omnis modi.", "Officiis perferendis iure sunt corporis iusto. Eveniet inventore autem accusamus neque placeat distinctio laborum. Voluptas voluptas et.", "Blanditiis nobis rerum quas et dolore. Mollitia dolorem quo voluptatibus eaque. Sapiente voluptatibus odit facere qui quos nostrum. Quos voluptatem ea voluptatem atque. Similique enim ex porro voluptas.", "Iusto debitis dolorum eius aperiam quibusdam. Molestias autem ut natus sequi quasi. Quam non aut voluptatem odio inventore dolores. Omnis ad vitae quia nostrum autem aut. Maxime rem consequatur."]