["Facere dignissimos facilis error qui voluptatem amet modi. Et velit pariatur voluptas est. Quia voluptate a sit qui quidem velit. Reiciendis temporibus error et itaque. Consequuntur debitis et doloremque sit quae maxime.", "Sint perferendis possimus tenetur numquam totam rerum. Laborum ipsa doloribus fugit debitis. Quibusdam voluptate dicta quidem et nemo ea magni. Quasi vel quod veniam sint eveniet. Aut sunt consectetur quia est recusandae ipsam in."]