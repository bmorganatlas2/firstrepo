["Dicta reprehenderit qui sed nulla unde natus. Odio aut qui at omnis libero. Mollitia nesciunt neque laudantium nisi sit.", "Quasi alias sapiente quibusdam quae. Quas iure exercitationem reiciendis et numquam velit. Ut quaerat inventore voluptate aperiam libero porro.", "Dolor ut deserunt nam quia vel autem. Fuga in tempora. Tenetur assumenda distinctio. Minus tempore sit. Consequatur ducimus occaecati.", "Quam omnis qui. Cupiditate aperiam eligendi voluptas. Nostrum unde iure culpa autem. Et sit quae quibusdam vero veritatis. Excepturi minima itaque possimus quas.", "Consequatur et sit vel. Est eius rerum nihil magni soluta officiis. Molestiae deleniti hic in rerum. Non architecto debitis laboriosam.", "Totam qui a consectetur nesciunt repellendus. Ea hic a debitis odio esse quo possimus. Rerum aut ipsam qui deleniti commodi dolore.", "Necessitatibus quia quo ullam. Earum quibusdam adipisci dicta est qui iste. Labore illum qui. Rerum asperiores aliquid et similique in iure. Fuga quod et adipisci pariatur velit sed inventore.", "Quos non et iure. Occaecati velit nobis quia expedita consequatur ducimus. Voluptatum est eos. Aperiam similique omnis.", "Tempora ut ea voluptatem magnam adipisci. Ut possimus repellendus eum reiciendis. Non occaecati sit aspernatur. Reiciendis ut totam ipsam aut veniam.", "Quis natus et. Soluta est dolorum aut maiores eos. Quis praesentium nulla et libero. Ipsam consectetur enim ipsa et harum est quis. Voluptatem et ut animi et cumque nobis ad."]