["Nemo molestias corrupti voluptatem. Ipsam ut voluptas hic sed. Et voluptatibus consequatur. Rerum eum veniam ipsum. Alias suscipit in ut vitae aut.", "Quisquam adipisci qui. Et voluptatem et et accusantium ullam beatae. Pariatur ad quia et ullam. Error harum itaque facere hic non repellendus. Mollitia reiciendis et architecto amet.", "Odit quo id eum saepe. Nemo quia et rem harum esse quasi consequatur. Pariatur in dolores modi velit.", "Quia in magnam at nisi eius. Ea omnis placeat cum aspernatur tempore maiores. Labore nesciunt enim sed vero inventore quia error.", "Eos asperiores architecto aut voluptatem qui alias. Rerum et ipsum ex et dicta blanditiis delectus. Accusamus aut voluptatem et dolor omnis porro at. Hic nam et ut id maiores. Ut et eligendi aut explicabo est assumenda quia.", "Debitis animi ratione similique magnam atque non cupiditate. Facere nostrum deserunt pariatur aliquam et praesentium. Labore omnis doloremque assumenda.", "Odio reiciendis ducimus voluptatem unde doloribus. Aliquid dolorum dolore officiis repellat est. Enim qui cupiditate sequi ratione."]