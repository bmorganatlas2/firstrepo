["Quo vitae fugiat error asperiores repellat ut delectus. In rerum ut sit rerum laudantium molestiae non. Asperiores voluptatem rerum excepturi. Ducimus provident et praesentium voluptatem in sint. Iusto quia ea.", "Est cumque fugiat aut cupiditate autem suscipit. Vel dolores ut molestiae a et provident perspiciatis. Perspiciatis voluptatem animi ab eligendi ipsam rerum maiores. Voluptatem aut at mollitia animi. Et voluptate minus aperiam et.", "Minima corrupti numquam autem. Rerum vero ab aperiam sint. Aut ullam impedit nihil at voluptatibus commodi.", "Rerum ut ab. Dolor perspiciatis harum repellendus. Non sint dolores recusandae. Facere omnis quibusdam ex consequatur. Aliquid tempora dicta consequatur aut excepturi.", "Et aut laborum. Sint magni enim officiis ut cum aperiam. Autem eius dolor amet ipsum ipsam. Tenetur molestias sunt quia quos est maiores. Vitae quam aut quas eum excepturi nesciunt quasi.", "Quas in eos voluptatem omnis est harum incidunt. Quod cum eum asperiores. Recusandae rem vitae odio et accusamus sint. Ratione id nihil id velit voluptatem. Minima labore impedit voluptatum ipsam eius."]