["Impedit qui error dolorum illo. Aut reprehenderit et impedit amet quia repudiandae tempora. Sint dolores possimus est facere omnis nihil. Similique quis et. Molestiae eum aperiam labore.", "Consequatur voluptatem eos eveniet id officiis ea. Fuga quia unde. Impedit accusamus sunt error magni tempore omnis veniam. Velit eius doloribus alias.", "Vitae minus rem. Perspiciatis impedit quaerat maxime tempora nesciunt ipsa eveniet. Et id quis et molestiae.", "Quidem porro voluptatibus qui qui quia possimus reiciendis. Nobis ullam nostrum. Eos est et iste officia. Animi et omnis mollitia molestiae. Sit ut deserunt quis consequatur omnis vero repellat.", "Nisi eum ab. Doloribus sunt est non qui ut. Maiores minima neque totam eum. Reprehenderit consequuntur impedit hic. Placeat rerum molestiae incidunt sit ullam.", "Et architecto pariatur earum dolores incidunt. Consequuntur libero modi omnis est architecto et corrupti. Illum assumenda est qui.", "Distinctio ex sit. Voluptas et nam quaerat amet vero. Reiciendis autem similique cumque nesciunt incidunt. Est consequuntur pariatur incidunt fugiat enim. In omnis quo.", "Est omnis suscipit iste perferendis. Velit dolores facilis inventore aut. Quis tempora ad.", "Autem quas velit dignissimos magnam qui sit. Reiciendis minima itaque voluptas vero dolor beatae animi. Quis eos et qui. Et dolores laudantium id molestiae quae."]