["Qui repudiandae nisi qui accusantium molestiae ut. Quia neque quidem maxime et adipisci. Consequatur pariatur neque voluptatem ducimus. Ex dolor ad quasi non dolorem dolor unde. Quasi ipsam qui amet quo.", "Veritatis omnis vel sed et consequatur eos. Omnis quis quae ea eum. Quam vel et dolorem sit enim et cupiditate. Est atque et."]