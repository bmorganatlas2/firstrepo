["Tempore animi provident laboriosam recusandae deserunt. Doloribus laboriosam aut est magni dignissimos aliquid et. Nesciunt voluptates quidem eius et possimus amet nemo. Saepe illum sit dignissimos dolor.", "Doloremque necessitatibus rem excepturi sunt in sit consectetur. Asperiores odit est. Vero quaerat consequatur odio cupiditate in quod sunt. Et impedit sapiente est nulla.", "Molestias et saepe. Exercitationem consequuntur at eos soluta ullam vero quaerat. Eum quos magnam temporibus. Sit repudiandae provident impedit quas. Esse voluptatibus illum quod suscipit nemo.", "Officiis quia est et recusandae quibusdam maxime molestiae. Nemo quia vel vitae facilis et aut nihil. Fugit necessitatibus aliquid quos. Vero nam cum corporis eaque ab. Est qui non omnis.", "Animi aperiam ea voluptas. Aut mollitia error. Est vel ullam rerum et.", "Eius qui eaque atque. Neque quo et quis voluptatem error. Sed saepe sit. Sed est expedita. Mollitia natus non rerum maxime.", "Tempore molestiae sed fuga voluptatem sint. Harum voluptatem sed dignissimos. In facere sequi et vitae commodi. Sunt nemo sapiente dolor rem inventore autem non.", "Voluptatibus iure est qui. Eligendi voluptas laborum asperiores sit eveniet. Temporibus eveniet aspernatur fuga. Ut voluptatum veritatis quas et. Rerum facilis voluptas quas vel omnis.", "Asperiores molestiae ducimus est. At nam est quia. Inventore ipsam consectetur sed id aperiam velit."]