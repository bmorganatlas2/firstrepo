["Sed quo qui rerum. Nihil unde fugiat sint nemo est. Totam qui quidem quaerat officia atque aliquid. Pariatur illum aliquid nihil quos.", "Quaerat culpa omnis et. Aspernatur ullam neque quia perferendis repellendus ex voluptas. Aut repudiandae tempore ut nulla ipsam ut.", "Non laboriosam qui est occaecati. Necessitatibus accusantium delectus dolorum voluptas aut. Voluptatem rem natus. Omnis magni corporis asperiores doloremque omnis voluptatem tempore.", "Atque cumque nisi quia quia ad aut. Totam et aut cum. Sint qui dolor. Dicta voluptate qui perferendis voluptatem laboriosam. Et harum itaque ut est sint ut enim.", "Aspernatur ad itaque. Sint reprehenderit ea sint corporis libero est veniam. Dolor perspiciatis assumenda architecto ex est sit. At maiores labore et molestiae. Autem sed itaque recusandae.", "Eius temporibus repellendus. Itaque alias magni officia tenetur quo adipisci. Molestiae repellat eos magni eligendi. Quas corrupti adipisci tempora. Necessitatibus autem deserunt culpa aut modi.", "Voluptas fuga aut animi velit quia laborum. Dignissimos ea voluptatem ab sint esse ut et. Eos rerum quia aspernatur. Hic quas commodi veniam recusandae quisquam id.", "Eius dolor sapiente fugiat. Iste eaque necessitatibus beatae. Nihil eos qui maxime non consectetur. Minima natus et quas suscipit nostrum. Nemo voluptatem assumenda officia a autem.", "Libero maxime quia quo repellendus qui nisi eum. Et nisi aut temporibus amet autem quia et. Rerum veritatis quia cumque laboriosam ut ipsum. Corrupti iure commodi vel consequatur illum totam."]