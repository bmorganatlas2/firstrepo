["Adipisci accusantium rerum. Quas aperiam quia laboriosam alias magni. Cupiditate qui eaque qui minus fugit voluptatem repudiandae.", "Suscipit quaerat iusto cupiditate voluptatem velit. Nihil autem recusandae rerum ipsam natus voluptate et. Id ullam a quod minima non. Mollitia est nobis est corporis.", "Adipisci ut rerum porro aut. Sint in perspiciatis omnis illo corporis quis. Et fugit voluptatem veritatis quia nihil fuga. Rerum numquam exercitationem qui deserunt nostrum aut accusantium. Dicta sed adipisci totam non deleniti.", "Delectus officiis ad vero. Laboriosam dignissimos minima quaerat qui eveniet omnis. Libero explicabo et aut distinctio accusantium mollitia. Non at maxime delectus corporis recusandae rem ipsum. Sed temporibus dolorum praesentium enim.", "Autem eos ad excepturi. Earum ducimus unde error consequatur sint quo occaecati. Debitis enim ex deleniti consequatur. Accusamus ea placeat officiis. Eveniet voluptas facilis nihil qui iure ut.", "Ut beatae voluptates vitae fugiat est illum. Deserunt nihil aperiam doloremque. Vel et nisi alias.", "Et quae earum facilis dicta officia aspernatur. Eum earum autem soluta. Iusto neque et nam et. Dolorem nihil tempora impedit inventore.", "Id alias iste qui in similique blanditiis. Voluptatem ipsum velit occaecati. Voluptatem libero veniam.", "Ad nulla voluptas nam. Incidunt sed sit consequuntur nisi ea nesciunt. Consequatur nihil eaque. Quaerat voluptas omnis inventore."]