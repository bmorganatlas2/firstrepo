["Similique dolor porro. Iste et excepturi asperiores ut. A eius quod et expedita libero quibusdam harum.", "Consequuntur non et et consequatur dolorum et mollitia. Ea dolores quam amet adipisci nostrum. Fugit praesentium nemo explicabo.", "Optio natus ratione. Eos illo recusandae. Odio fuga repellendus modi enim sit. Laborum aliquam aut consectetur nam est totam. Deleniti neque sint quae et ut eos mollitia."]